netcdf trentino_hourlyweatherdata {
dimensions:
	Station = UNLIMITED ; // (3 currently)
	characters = 200 ;
	Time = UNLIMITED ; // (17520 currently)
variables:
	int Station(Station) ;
		Station:units = "id" ;
		Station:long_name = "Station" ;
	double StationLat(Station) ;
		StationLat:units = "degrees North" ;
		StationLat:_FillValue = NaN ;
	double StationLon(Station) ;
		StationLon:units = "degrees East" ;
		StationLon:_FillValue = NaN ;
	char StationIdName(Station, characters) ;
	double Time(Time) ;
		Time:units = "senconds since 1970-01-01 +1" ;
		Time:long_name = "Time" ;
	double Prec(Time, Station) ;
		Prec:units = "millimeters" ;
		Prec:_FillValue = NaN ;
		Prec:long_name = "Hourly Precipitation" ;
	double Temp(Time, Station) ;
		Temp:units = "degrees C" ;
		Temp:_FillValue = NaN ;
		Temp:long_name = "Averaged Air Temperature" ;
data:

 Station = 1, 2, 3 ;

 StationLat = 45.886196, 46.194763, 46.014465 ;

 StationLon = 10.944168, 11.169777, 10.866802 ;

 StationIdName =
  "FEMst21",
  "FEMst22",
  "FEMst23" ;

 Time = 1109635200, 1109638800, 1109642400, 1109646000, 1109649600, 
    1109653200, 1109656800, 1109660400, 1109664000, 1109667600, 1109671200, 
    1109674800, 1109678400, 1109682000, 1109685600, 1109689200, 1109692800, 
    1109696400, 1109700000, 1109703600, 1109707200, 1109710800, 1109714400, 
    1109718000, 1109721600, 1109725200, 1109728800, 1109732400, 1109736000, 
    1109739600, 1109743200, 1109746800, 1109750400, 1109754000, 1109757600, 
    1109761200, 1109764800, 1109768400, 1109772000, 1109775600, 1109779200, 
    1109782800, 1109786400, 1109790000, 1109793600, 1109797200, 1109800800, 
    1109804400, 1109808000, 1109811600, 1109815200, 1109818800, 1109822400, 
    1109826000, 1109829600, 1109833200, 1109836800, 1109840400, 1109844000, 
    1109847600, 1109851200, 1109854800, 1109858400, 1109862000, 1109865600, 
    1109869200, 1109872800, 1109876400, 1109880000, 1109883600, 1109887200, 
    1109890800, 1109894400, 1109898000, 1109901600, 1109905200, 1109908800, 
    1109912400, 1109916000, 1109919600, 1109923200, 1109926800, 1109930400, 
    1109934000, 1109937600, 1109941200, 1109944800, 1109948400, 1109952000, 
    1109955600, 1109959200, 1109962800, 1109966400, 1109970000, 1109973600, 
    1109977200, 1109980800, 1109984400, 1109988000, 1109991600, 1109995200, 
    1109998800, 1110002400, 1110006000, 1110009600, 1110013200, 1110016800, 
    1110020400, 1110024000, 1110027600, 1110031200, 1110034800, 1110038400, 
    1110042000, 1110045600, 1110049200, 1110052800, 1110056400, 1110060000, 
    1110063600, 1110067200, 1110070800, 1110074400, 1110078000, 1110081600, 
    1110085200, 1110088800, 1110092400, 1110096000, 1110099600, 1110103200, 
    1110106800, 1110110400, 1110114000, 1110117600, 1110121200, 1110124800, 
    1110128400, 1110132000, 1110135600, 1110139200, 1110142800, 1110146400, 
    1110150000, 1110153600, 1110157200, 1110160800, 1110164400, 1110168000, 
    1110171600, 1110175200, 1110178800, 1110182400, 1110186000, 1110189600, 
    1110193200, 1110196800, 1110200400, 1110204000, 1110207600, 1110211200, 
    1110214800, 1110218400, 1110222000, 1110225600, 1110229200, 1110232800, 
    1110236400, 1110240000, 1110243600, 1110247200, 1110250800, 1110254400, 
    1110258000, 1110261600, 1110265200, 1110268800, 1110272400, 1110276000, 
    1110279600, 1110283200, 1110286800, 1110290400, 1110294000, 1110297600, 
    1110301200, 1110304800, 1110308400, 1110312000, 1110315600, 1110319200, 
    1110322800, 1110326400, 1110330000, 1110333600, 1110337200, 1110340800, 
    1110344400, 1110348000, 1110351600, 1110355200, 1110358800, 1110362400, 
    1110366000, 1110369600, 1110373200, 1110376800, 1110380400, 1110384000, 
    1110387600, 1110391200, 1110394800, 1110398400, 1110402000, 1110405600, 
    1110409200, 1110412800, 1110416400, 1110420000, 1110423600, 1110427200, 
    1110430800, 1110434400, 1110438000, 1110441600, 1110445200, 1110448800, 
    1110452400, 1110456000, 1110459600, 1110463200, 1110466800, 1110470400, 
    1110474000, 1110477600, 1110481200, 1110484800, 1110488400, 1110492000, 
    1110495600, 1110499200, 1110502800, 1110506400, 1110510000, 1110513600, 
    1110517200, 1110520800, 1110524400, 1110528000, 1110531600, 1110535200, 
    1110538800, 1110542400, 1110546000, 1110549600, 1110553200, 1110556800, 
    1110560400, 1110564000, 1110567600, 1110571200, 1110574800, 1110578400, 
    1110582000, 1110585600, 1110589200, 1110592800, 1110596400, 1110600000, 
    1110603600, 1110607200, 1110610800, 1110614400, 1110618000, 1110621600, 
    1110625200, 1110628800, 1110632400, 1110636000, 1110639600, 1110643200, 
    1110646800, 1110650400, 1110654000, 1110657600, 1110661200, 1110664800, 
    1110668400, 1110672000, 1110675600, 1110679200, 1110682800, 1110686400, 
    1110690000, 1110693600, 1110697200, 1110700800, 1110704400, 1110708000, 
    1110711600, 1110715200, 1110718800, 1110722400, 1110726000, 1110729600, 
    1110733200, 1110736800, 1110740400, 1110744000, 1110747600, 1110751200, 
    1110754800, 1110758400, 1110762000, 1110765600, 1110769200, 1110772800, 
    1110776400, 1110780000, 1110783600, 1110787200, 1110790800, 1110794400, 
    1110798000, 1110801600, 1110805200, 1110808800, 1110812400, 1110816000, 
    1110819600, 1110823200, 1110826800, 1110830400, 1110834000, 1110837600, 
    1110841200, 1110844800, 1110848400, 1110852000, 1110855600, 1110859200, 
    1110862800, 1110866400, 1110870000, 1110873600, 1110877200, 1110880800, 
    1110884400, 1110888000, 1110891600, 1110895200, 1110898800, 1110902400, 
    1110906000, 1110909600, 1110913200, 1110916800, 1110920400, 1110924000, 
    1110927600, 1110931200, 1110934800, 1110938400, 1110942000, 1110945600, 
    1110949200, 1110952800, 1110956400, 1110960000, 1110963600, 1110967200, 
    1110970800, 1110974400, 1110978000, 1110981600, 1110985200, 1110988800, 
    1110992400, 1110996000, 1110999600, 1111003200, 1111006800, 1111010400, 
    1111014000, 1111017600, 1111021200, 1111024800, 1111028400, 1111032000, 
    1111035600, 1111039200, 1111042800, 1111046400, 1111050000, 1111053600, 
    1111057200, 1111060800, 1111064400, 1111068000, 1111071600, 1111075200, 
    1111078800, 1111082400, 1111086000, 1111089600, 1111093200, 1111096800, 
    1111100400, 1111104000, 1111107600, 1111111200, 1111114800, 1111118400, 
    1111122000, 1111125600, 1111129200, 1111132800, 1111136400, 1111140000, 
    1111143600, 1111147200, 1111150800, 1111154400, 1111158000, 1111161600, 
    1111165200, 1111168800, 1111172400, 1111176000, 1111179600, 1111183200, 
    1111186800, 1111190400, 1111194000, 1111197600, 1111201200, 1111204800, 
    1111208400, 1111212000, 1111215600, 1111219200, 1111222800, 1111226400, 
    1111230000, 1111233600, 1111237200, 1111240800, 1111244400, 1111248000, 
    1111251600, 1111255200, 1111258800, 1111262400, 1111266000, 1111269600, 
    1111273200, 1111276800, 1111280400, 1111284000, 1111287600, 1111291200, 
    1111294800, 1111298400, 1111302000, 1111305600, 1111309200, 1111312800, 
    1111316400, 1111320000, 1111323600, 1111327200, 1111330800, 1111334400, 
    1111338000, 1111341600, 1111345200, 1111348800, 1111352400, 1111356000, 
    1111359600, 1111363200, 1111366800, 1111370400, 1111374000, 1111377600, 
    1111381200, 1111384800, 1111388400, 1111392000, 1111395600, 1111399200, 
    1111402800, 1111406400, 1111410000, 1111413600, 1111417200, 1111420800, 
    1111424400, 1111428000, 1111431600, 1111435200, 1111438800, 1111442400, 
    1111446000, 1111449600, 1111453200, 1111456800, 1111460400, 1111464000, 
    1111467600, 1111471200, 1111474800, 1111478400, 1111482000, 1111485600, 
    1111489200, 1111492800, 1111496400, 1111500000, 1111503600, 1111507200, 
    1111510800, 1111514400, 1111518000, 1111521600, 1111525200, 1111528800, 
    1111532400, 1111536000, 1111539600, 1111543200, 1111546800, 1111550400, 
    1111554000, 1111557600, 1111561200, 1111564800, 1111568400, 1111572000, 
    1111575600, 1111579200, 1111582800, 1111586400, 1111590000, 1111593600, 
    1111597200, 1111600800, 1111604400, 1111608000, 1111611600, 1111615200, 
    1111618800, 1111622400, 1111626000, 1111629600, 1111633200, 1111636800, 
    1111640400, 1111644000, 1111647600, 1111651200, 1111654800, 1111658400, 
    1111662000, 1111665600, 1111669200, 1111672800, 1111676400, 1111680000, 
    1111683600, 1111687200, 1111690800, 1111694400, 1111698000, 1111701600, 
    1111705200, 1111708800, 1111712400, 1111716000, 1111719600, 1111723200, 
    1111726800, 1111730400, 1111734000, 1111737600, 1111741200, 1111744800, 
    1111748400, 1111752000, 1111755600, 1111759200, 1111762800, 1111766400, 
    1111770000, 1111773600, 1111777200, 1111780800, 1111784400, 1111788000, 
    1111791600, 1111795200, 1111798800, 1111802400, 1111806000, 1111809600, 
    1111813200, 1111816800, 1111820400, 1111824000, 1111827600, 1111831200, 
    1111834800, 1111838400, 1111842000, 1111845600, 1111849200, 1111852800, 
    1111856400, 1111860000, 1111863600, 1111867200, 1111870800, 1111874400, 
    1111878000, 1111881600, 1111885200, 1111888800, 1111892400, 1111896000, 
    1111899600, 1111903200, 1111906800, 1111910400, 1111914000, 1111917600, 
    1111921200, 1111924800, 1111928400, 1111932000, 1111935600, 1111939200, 
    1111942800, 1111946400, 1111950000, 1111953600, 1111957200, 1111960800, 
    1111964400, 1111968000, 1111971600, 1111975200, 1111978800, 1111982400, 
    1111986000, 1111989600, 1111993200, 1111996800, 1112000400, 1112004000, 
    1112007600, 1112011200, 1112014800, 1112018400, 1112022000, 1112025600, 
    1112029200, 1112032800, 1112036400, 1112040000, 1112043600, 1112047200, 
    1112050800, 1112054400, 1112058000, 1112061600, 1112065200, 1112068800, 
    1112072400, 1112076000, 1112079600, 1112083200, 1112086800, 1112090400, 
    1112094000, 1112097600, 1112101200, 1112104800, 1112108400, 1112112000, 
    1112115600, 1112119200, 1112122800, 1112126400, 1112130000, 1112133600, 
    1112137200, 1112140800, 1112144400, 1112148000, 1112151600, 1112155200, 
    1112158800, 1112162400, 1112166000, 1112169600, 1112173200, 1112176800, 
    1112180400, 1112184000, 1112187600, 1112191200, 1112194800, 1112198400, 
    1112202000, 1112205600, 1112209200, 1112212800, 1112216400, 1112220000, 
    1112223600, 1112227200, 1112230800, 1112234400, 1112238000, 1112241600, 
    1112245200, 1112248800, 1112252400, 1112256000, 1112259600, 1112263200, 
    1112266800, 1112270400, 1112274000, 1112277600, 1112281200, 1112284800, 
    1112288400, 1112292000, 1112295600, 1112299200, 1112302800, 1112306400, 
    1112310000, 1112313600, 1112317200, 1112320800, 1112324400, 1112328000, 
    1112331600, 1112335200, 1112338800, 1112342400, 1112346000, 1112349600, 
    1112353200, 1112356800, 1112360400, 1112364000, 1112367600, 1112371200, 
    1112374800, 1112378400, 1112382000, 1112385600, 1112389200, 1112392800, 
    1112396400, 1112400000, 1112403600, 1112407200, 1112410800, 1112414400, 
    1112418000, 1112421600, 1112425200, 1112428800, 1112432400, 1112436000, 
    1112439600, 1112443200, 1112446800, 1112450400, 1112454000, 1112457600, 
    1112461200, 1112464800, 1112468400, 1112472000, 1112475600, 1112479200, 
    1112482800, 1112486400, 1112490000, 1112493600, 1112497200, 1112500800, 
    1112504400, 1112508000, 1112511600, 1112515200, 1112518800, 1112522400, 
    1112526000, 1112529600, 1112533200, 1112536800, 1112540400, 1112544000, 
    1112547600, 1112551200, 1112554800, 1112558400, 1112562000, 1112565600, 
    1112569200, 1112572800, 1112576400, 1112580000, 1112583600, 1112587200, 
    1112590800, 1112594400, 1112598000, 1112601600, 1112605200, 1112608800, 
    1112612400, 1112616000, 1112619600, 1112623200, 1112626800, 1112630400, 
    1112634000, 1112637600, 1112641200, 1112644800, 1112648400, 1112652000, 
    1112655600, 1112659200, 1112662800, 1112666400, 1112670000, 1112673600, 
    1112677200, 1112680800, 1112684400, 1112688000, 1112691600, 1112695200, 
    1112698800, 1112702400, 1112706000, 1112709600, 1112713200, 1112716800, 
    1112720400, 1112724000, 1112727600, 1112731200, 1112734800, 1112738400, 
    1112742000, 1112745600, 1112749200, 1112752800, 1112756400, 1112760000, 
    1112763600, 1112767200, 1112770800, 1112774400, 1112778000, 1112781600, 
    1112785200, 1112788800, 1112792400, 1112796000, 1112799600, 1112803200, 
    1112806800, 1112810400, 1112814000, 1112817600, 1112821200, 1112824800, 
    1112828400, 1112832000, 1112835600, 1112839200, 1112842800, 1112846400, 
    1112850000, 1112853600, 1112857200, 1112860800, 1112864400, 1112868000, 
    1112871600, 1112875200, 1112878800, 1112882400, 1112886000, 1112889600, 
    1112893200, 1112896800, 1112900400, 1112904000, 1112907600, 1112911200, 
    1112914800, 1112918400, 1112922000, 1112925600, 1112929200, 1112932800, 
    1112936400, 1112940000, 1112943600, 1112947200, 1112950800, 1112954400, 
    1112958000, 1112961600, 1112965200, 1112968800, 1112972400, 1112976000, 
    1112979600, 1112983200, 1112986800, 1112990400, 1112994000, 1112997600, 
    1113001200, 1113004800, 1113008400, 1113012000, 1113015600, 1113019200, 
    1113022800, 1113026400, 1113030000, 1113033600, 1113037200, 1113040800, 
    1113044400, 1113048000, 1113051600, 1113055200, 1113058800, 1113062400, 
    1113066000, 1113069600, 1113073200, 1113076800, 1113080400, 1113084000, 
    1113087600, 1113091200, 1113094800, 1113098400, 1113102000, 1113105600, 
    1113109200, 1113112800, 1113116400, 1113120000, 1113123600, 1113127200, 
    1113130800, 1113134400, 1113138000, 1113141600, 1113145200, 1113148800, 
    1113152400, 1113156000, 1113159600, 1113163200, 1113166800, 1113170400, 
    1113174000, 1113177600, 1113181200, 1113184800, 1113188400, 1113192000, 
    1113195600, 1113199200, 1113202800, 1113206400, 1113210000, 1113213600, 
    1113217200, 1113220800, 1113224400, 1113228000, 1113231600, 1113235200, 
    1113238800, 1113242400, 1113246000, 1113249600, 1113253200, 1113256800, 
    1113260400, 1113264000, 1113267600, 1113271200, 1113274800, 1113278400, 
    1113282000, 1113285600, 1113289200, 1113292800, 1113296400, 1113300000, 
    1113303600, 1113307200, 1113310800, 1113314400, 1113318000, 1113321600, 
    1113325200, 1113328800, 1113332400, 1113336000, 1113339600, 1113343200, 
    1113346800, 1113350400, 1113354000, 1113357600, 1113361200, 1113364800, 
    1113368400, 1113372000, 1113375600, 1113379200, 1113382800, 1113386400, 
    1113390000, 1113393600, 1113397200, 1113400800, 1113404400, 1113408000, 
    1113411600, 1113415200, 1113418800, 1113422400, 1113426000, 1113429600, 
    1113433200, 1113436800, 1113440400, 1113444000, 1113447600, 1113451200, 
    1113454800, 1113458400, 1113462000, 1113465600, 1113469200, 1113472800, 
    1113476400, 1113480000, 1113483600, 1113487200, 1113490800, 1113494400, 
    1113498000, 1113501600, 1113505200, 1113508800, 1113512400, 1113516000, 
    1113519600, 1113523200, 1113526800, 1113530400, 1113534000, 1113537600, 
    1113541200, 1113544800, 1113548400, 1113552000, 1113555600, 1113559200, 
    1113562800, 1113566400, 1113570000, 1113573600, 1113577200, 1113580800, 
    1113584400, 1113588000, 1113591600, 1113595200, 1113598800, 1113602400, 
    1113606000, 1113609600, 1113613200, 1113616800, 1113620400, 1113624000, 
    1113627600, 1113631200, 1113634800, 1113638400, 1113642000, 1113645600, 
    1113649200, 1113652800, 1113656400, 1113660000, 1113663600, 1113667200, 
    1113670800, 1113674400, 1113678000, 1113681600, 1113685200, 1113688800, 
    1113692400, 1113696000, 1113699600, 1113703200, 1113706800, 1113710400, 
    1113714000, 1113717600, 1113721200, 1113724800, 1113728400, 1113732000, 
    1113735600, 1113739200, 1113742800, 1113746400, 1113750000, 1113753600, 
    1113757200, 1113760800, 1113764400, 1113768000, 1113771600, 1113775200, 
    1113778800, 1113782400, 1113786000, 1113789600, 1113793200, 1113796800, 
    1113800400, 1113804000, 1113807600, 1113811200, 1113814800, 1113818400, 
    1113822000, 1113825600, 1113829200, 1113832800, 1113836400, 1113840000, 
    1113843600, 1113847200, 1113850800, 1113854400, 1113858000, 1113861600, 
    1113865200, 1113868800, 1113872400, 1113876000, 1113879600, 1113883200, 
    1113886800, 1113890400, 1113894000, 1113897600, 1113901200, 1113904800, 
    1113908400, 1113912000, 1113915600, 1113919200, 1113922800, 1113926400, 
    1113930000, 1113933600, 1113937200, 1113940800, 1113944400, 1113948000, 
    1113951600, 1113955200, 1113958800, 1113962400, 1113966000, 1113969600, 
    1113973200, 1113976800, 1113980400, 1113984000, 1113987600, 1113991200, 
    1113994800, 1113998400, 1114002000, 1114005600, 1114009200, 1114012800, 
    1114016400, 1114020000, 1114023600, 1114027200, 1114030800, 1114034400, 
    1114038000, 1114041600, 1114045200, 1114048800, 1114052400, 1114056000, 
    1114059600, 1114063200, 1114066800, 1114070400, 1114074000, 1114077600, 
    1114081200, 1114084800, 1114088400, 1114092000, 1114095600, 1114099200, 
    1114102800, 1114106400, 1114110000, 1114113600, 1114117200, 1114120800, 
    1114124400, 1114128000, 1114131600, 1114135200, 1114138800, 1114142400, 
    1114146000, 1114149600, 1114153200, 1114156800, 1114160400, 1114164000, 
    1114167600, 1114171200, 1114174800, 1114178400, 1114182000, 1114185600, 
    1114189200, 1114192800, 1114196400, 1114200000, 1114203600, 1114207200, 
    1114210800, 1114214400, 1114218000, 1114221600, 1114225200, 1114228800, 
    1114232400, 1114236000, 1114239600, 1114243200, 1114246800, 1114250400, 
    1114254000, 1114257600, 1114261200, 1114264800, 1114268400, 1114272000, 
    1114275600, 1114279200, 1114282800, 1114286400, 1114290000, 1114293600, 
    1114297200, 1114300800, 1114304400, 1114308000, 1114311600, 1114315200, 
    1114318800, 1114322400, 1114326000, 1114329600, 1114333200, 1114336800, 
    1114340400, 1114344000, 1114347600, 1114351200, 1114354800, 1114358400, 
    1114362000, 1114365600, 1114369200, 1114372800, 1114376400, 1114380000, 
    1114383600, 1114387200, 1114390800, 1114394400, 1114398000, 1114401600, 
    1114405200, 1114408800, 1114412400, 1114416000, 1114419600, 1114423200, 
    1114426800, 1114430400, 1114434000, 1114437600, 1114441200, 1114444800, 
    1114448400, 1114452000, 1114455600, 1114459200, 1114462800, 1114466400, 
    1114470000, 1114473600, 1114477200, 1114480800, 1114484400, 1114488000, 
    1114491600, 1114495200, 1114498800, 1114502400, 1114506000, 1114509600, 
    1114513200, 1114516800, 1114520400, 1114524000, 1114527600, 1114531200, 
    1114534800, 1114538400, 1114542000, 1114545600, 1114549200, 1114552800, 
    1114556400, 1114560000, 1114563600, 1114567200, 1114570800, 1114574400, 
    1114578000, 1114581600, 1114585200, 1114588800, 1114592400, 1114596000, 
    1114599600, 1114603200, 1114606800, 1114610400, 1114614000, 1114617600, 
    1114621200, 1114624800, 1114628400, 1114632000, 1114635600, 1114639200, 
    1114642800, 1114646400, 1114650000, 1114653600, 1114657200, 1114660800, 
    1114664400, 1114668000, 1114671600, 1114675200, 1114678800, 1114682400, 
    1114686000, 1114689600, 1114693200, 1114696800, 1114700400, 1114704000, 
    1114707600, 1114711200, 1114714800, 1114718400, 1114722000, 1114725600, 
    1114729200, 1114732800, 1114736400, 1114740000, 1114743600, 1114747200, 
    1114750800, 1114754400, 1114758000, 1114761600, 1114765200, 1114768800, 
    1114772400, 1114776000, 1114779600, 1114783200, 1114786800, 1114790400, 
    1114794000, 1114797600, 1114801200, 1114804800, 1114808400, 1114812000, 
    1114815600, 1114819200, 1114822800, 1114826400, 1114830000, 1114833600, 
    1114837200, 1114840800, 1114844400, 1114848000, 1114851600, 1114855200, 
    1114858800, 1114862400, 1114866000, 1114869600, 1114873200, 1114876800, 
    1114880400, 1114884000, 1114887600, 1114891200, 1114894800, 1114898400, 
    1114902000, 1114905600, 1114909200, 1114912800, 1114916400, 1114920000, 
    1114923600, 1114927200, 1114930800, 1114934400, 1114938000, 1114941600, 
    1114945200, 1114948800, 1114952400, 1114956000, 1114959600, 1114963200, 
    1114966800, 1114970400, 1114974000, 1114977600, 1114981200, 1114984800, 
    1114988400, 1114992000, 1114995600, 1114999200, 1115002800, 1115006400, 
    1115010000, 1115013600, 1115017200, 1115020800, 1115024400, 1115028000, 
    1115031600, 1115035200, 1115038800, 1115042400, 1115046000, 1115049600, 
    1115053200, 1115056800, 1115060400, 1115064000, 1115067600, 1115071200, 
    1115074800, 1115078400, 1115082000, 1115085600, 1115089200, 1115092800, 
    1115096400, 1115100000, 1115103600, 1115107200, 1115110800, 1115114400, 
    1115118000, 1115121600, 1115125200, 1115128800, 1115132400, 1115136000, 
    1115139600, 1115143200, 1115146800, 1115150400, 1115154000, 1115157600, 
    1115161200, 1115164800, 1115168400, 1115172000, 1115175600, 1115179200, 
    1115182800, 1115186400, 1115190000, 1115193600, 1115197200, 1115200800, 
    1115204400, 1115208000, 1115211600, 1115215200, 1115218800, 1115222400, 
    1115226000, 1115229600, 1115233200, 1115236800, 1115240400, 1115244000, 
    1115247600, 1115251200, 1115254800, 1115258400, 1115262000, 1115265600, 
    1115269200, 1115272800, 1115276400, 1115280000, 1115283600, 1115287200, 
    1115290800, 1115294400, 1115298000, 1115301600, 1115305200, 1115308800, 
    1115312400, 1115316000, 1115319600, 1115323200, 1115326800, 1115330400, 
    1115334000, 1115337600, 1115341200, 1115344800, 1115348400, 1115352000, 
    1115355600, 1115359200, 1115362800, 1115366400, 1115370000, 1115373600, 
    1115377200, 1115380800, 1115384400, 1115388000, 1115391600, 1115395200, 
    1115398800, 1115402400, 1115406000, 1115409600, 1115413200, 1115416800, 
    1115420400, 1115424000, 1115427600, 1115431200, 1115434800, 1115438400, 
    1115442000, 1115445600, 1115449200, 1115452800, 1115456400, 1115460000, 
    1115463600, 1115467200, 1115470800, 1115474400, 1115478000, 1115481600, 
    1115485200, 1115488800, 1115492400, 1115496000, 1115499600, 1115503200, 
    1115506800, 1115510400, 1115514000, 1115517600, 1115521200, 1115524800, 
    1115528400, 1115532000, 1115535600, 1115539200, 1115542800, 1115546400, 
    1115550000, 1115553600, 1115557200, 1115560800, 1115564400, 1115568000, 
    1115571600, 1115575200, 1115578800, 1115582400, 1115586000, 1115589600, 
    1115593200, 1115596800, 1115600400, 1115604000, 1115607600, 1115611200, 
    1115614800, 1115618400, 1115622000, 1115625600, 1115629200, 1115632800, 
    1115636400, 1115640000, 1115643600, 1115647200, 1115650800, 1115654400, 
    1115658000, 1115661600, 1115665200, 1115668800, 1115672400, 1115676000, 
    1115679600, 1115683200, 1115686800, 1115690400, 1115694000, 1115697600, 
    1115701200, 1115704800, 1115708400, 1115712000, 1115715600, 1115719200, 
    1115722800, 1115726400, 1115730000, 1115733600, 1115737200, 1115740800, 
    1115744400, 1115748000, 1115751600, 1115755200, 1115758800, 1115762400, 
    1115766000, 1115769600, 1115773200, 1115776800, 1115780400, 1115784000, 
    1115787600, 1115791200, 1115794800, 1115798400, 1115802000, 1115805600, 
    1115809200, 1115812800, 1115816400, 1115820000, 1115823600, 1115827200, 
    1115830800, 1115834400, 1115838000, 1115841600, 1115845200, 1115848800, 
    1115852400, 1115856000, 1115859600, 1115863200, 1115866800, 1115870400, 
    1115874000, 1115877600, 1115881200, 1115884800, 1115888400, 1115892000, 
    1115895600, 1115899200, 1115902800, 1115906400, 1115910000, 1115913600, 
    1115917200, 1115920800, 1115924400, 1115928000, 1115931600, 1115935200, 
    1115938800, 1115942400, 1115946000, 1115949600, 1115953200, 1115956800, 
    1115960400, 1115964000, 1115967600, 1115971200, 1115974800, 1115978400, 
    1115982000, 1115985600, 1115989200, 1115992800, 1115996400, 1116000000, 
    1116003600, 1116007200, 1116010800, 1116014400, 1116018000, 1116021600, 
    1116025200, 1116028800, 1116032400, 1116036000, 1116039600, 1116043200, 
    1116046800, 1116050400, 1116054000, 1116057600, 1116061200, 1116064800, 
    1116068400, 1116072000, 1116075600, 1116079200, 1116082800, 1116086400, 
    1116090000, 1116093600, 1116097200, 1116100800, 1116104400, 1116108000, 
    1116111600, 1116115200, 1116118800, 1116122400, 1116126000, 1116129600, 
    1116133200, 1116136800, 1116140400, 1116144000, 1116147600, 1116151200, 
    1116154800, 1116158400, 1116162000, 1116165600, 1116169200, 1116172800, 
    1116176400, 1116180000, 1116183600, 1116187200, 1116190800, 1116194400, 
    1116198000, 1116201600, 1116205200, 1116208800, 1116212400, 1116216000, 
    1116219600, 1116223200, 1116226800, 1116230400, 1116234000, 1116237600, 
    1116241200, 1116244800, 1116248400, 1116252000, 1116255600, 1116259200, 
    1116262800, 1116266400, 1116270000, 1116273600, 1116277200, 1116280800, 
    1116284400, 1116288000, 1116291600, 1116295200, 1116298800, 1116302400, 
    1116306000, 1116309600, 1116313200, 1116316800, 1116320400, 1116324000, 
    1116327600, 1116331200, 1116334800, 1116338400, 1116342000, 1116345600, 
    1116349200, 1116352800, 1116356400, 1116360000, 1116363600, 1116367200, 
    1116370800, 1116374400, 1116378000, 1116381600, 1116385200, 1116388800, 
    1116392400, 1116396000, 1116399600, 1116403200, 1116406800, 1116410400, 
    1116414000, 1116417600, 1116421200, 1116424800, 1116428400, 1116432000, 
    1116435600, 1116439200, 1116442800, 1116446400, 1116450000, 1116453600, 
    1116457200, 1116460800, 1116464400, 1116468000, 1116471600, 1116475200, 
    1116478800, 1116482400, 1116486000, 1116489600, 1116493200, 1116496800, 
    1116500400, 1116504000, 1116507600, 1116511200, 1116514800, 1116518400, 
    1116522000, 1116525600, 1116529200, 1116532800, 1116536400, 1116540000, 
    1116543600, 1116547200, 1116550800, 1116554400, 1116558000, 1116561600, 
    1116565200, 1116568800, 1116572400, 1116576000, 1116579600, 1116583200, 
    1116586800, 1116590400, 1116594000, 1116597600, 1116601200, 1116604800, 
    1116608400, 1116612000, 1116615600, 1116619200, 1116622800, 1116626400, 
    1116630000, 1116633600, 1116637200, 1116640800, 1116644400, 1116648000, 
    1116651600, 1116655200, 1116658800, 1116662400, 1116666000, 1116669600, 
    1116673200, 1116676800, 1116680400, 1116684000, 1116687600, 1116691200, 
    1116694800, 1116698400, 1116702000, 1116705600, 1116709200, 1116712800, 
    1116716400, 1116720000, 1116723600, 1116727200, 1116730800, 1116734400, 
    1116738000, 1116741600, 1116745200, 1116748800, 1116752400, 1116756000, 
    1116759600, 1116763200, 1116766800, 1116770400, 1116774000, 1116777600, 
    1116781200, 1116784800, 1116788400, 1116792000, 1116795600, 1116799200, 
    1116802800, 1116806400, 1116810000, 1116813600, 1116817200, 1116820800, 
    1116824400, 1116828000, 1116831600, 1116835200, 1116838800, 1116842400, 
    1116846000, 1116849600, 1116853200, 1116856800, 1116860400, 1116864000, 
    1116867600, 1116871200, 1116874800, 1116878400, 1116882000, 1116885600, 
    1116889200, 1116892800, 1116896400, 1116900000, 1116903600, 1116907200, 
    1116910800, 1116914400, 1116918000, 1116921600, 1116925200, 1116928800, 
    1116932400, 1116936000, 1116939600, 1116943200, 1116946800, 1116950400, 
    1116954000, 1116957600, 1116961200, 1116964800, 1116968400, 1116972000, 
    1116975600, 1116979200, 1116982800, 1116986400, 1116990000, 1116993600, 
    1116997200, 1117000800, 1117004400, 1117008000, 1117011600, 1117015200, 
    1117018800, 1117022400, 1117026000, 1117029600, 1117033200, 1117036800, 
    1117040400, 1117044000, 1117047600, 1117051200, 1117054800, 1117058400, 
    1117062000, 1117065600, 1117069200, 1117072800, 1117076400, 1117080000, 
    1117083600, 1117087200, 1117090800, 1117094400, 1117098000, 1117101600, 
    1117105200, 1117108800, 1117112400, 1117116000, 1117119600, 1117123200, 
    1117126800, 1117130400, 1117134000, 1117137600, 1117141200, 1117144800, 
    1117148400, 1117152000, 1117155600, 1117159200, 1117162800, 1117166400, 
    1117170000, 1117173600, 1117177200, 1117180800, 1117184400, 1117188000, 
    1117191600, 1117195200, 1117198800, 1117202400, 1117206000, 1117209600, 
    1117213200, 1117216800, 1117220400, 1117224000, 1117227600, 1117231200, 
    1117234800, 1117238400, 1117242000, 1117245600, 1117249200, 1117252800, 
    1117256400, 1117260000, 1117263600, 1117267200, 1117270800, 1117274400, 
    1117278000, 1117281600, 1117285200, 1117288800, 1117292400, 1117296000, 
    1117299600, 1117303200, 1117306800, 1117310400, 1117314000, 1117317600, 
    1117321200, 1117324800, 1117328400, 1117332000, 1117335600, 1117339200, 
    1117342800, 1117346400, 1117350000, 1117353600, 1117357200, 1117360800, 
    1117364400, 1117368000, 1117371600, 1117375200, 1117378800, 1117382400, 
    1117386000, 1117389600, 1117393200, 1117396800, 1117400400, 1117404000, 
    1117407600, 1117411200, 1117414800, 1117418400, 1117422000, 1117425600, 
    1117429200, 1117432800, 1117436400, 1117440000, 1117443600, 1117447200, 
    1117450800, 1117454400, 1117458000, 1117461600, 1117465200, 1117468800, 
    1117472400, 1117476000, 1117479600, 1117483200, 1117486800, 1117490400, 
    1117494000, 1117497600, 1117501200, 1117504800, 1117508400, 1117512000, 
    1117515600, 1117519200, 1117522800, 1117526400, 1117530000, 1117533600, 
    1117537200, 1117540800, 1117544400, 1117548000, 1117551600, 1117555200, 
    1117558800, 1117562400, 1117566000, 1117569600, 1117573200, 1117576800, 
    1117580400, 1117584000, 1117587600, 1117591200, 1117594800, 1117598400, 
    1117602000, 1117605600, 1117609200, 1117612800, 1117616400, 1117620000, 
    1117623600, 1117627200, 1117630800, 1117634400, 1117638000, 1117641600, 
    1117645200, 1117648800, 1117652400, 1117656000, 1117659600, 1117663200, 
    1117666800, 1117670400, 1117674000, 1117677600, 1117681200, 1117684800, 
    1117688400, 1117692000, 1117695600, 1117699200, 1117702800, 1117706400, 
    1117710000, 1117713600, 1117717200, 1117720800, 1117724400, 1117728000, 
    1117731600, 1117735200, 1117738800, 1117742400, 1117746000, 1117749600, 
    1117753200, 1117756800, 1117760400, 1117764000, 1117767600, 1117771200, 
    1117774800, 1117778400, 1117782000, 1117785600, 1117789200, 1117792800, 
    1117796400, 1117800000, 1117803600, 1117807200, 1117810800, 1117814400, 
    1117818000, 1117821600, 1117825200, 1117828800, 1117832400, 1117836000, 
    1117839600, 1117843200, 1117846800, 1117850400, 1117854000, 1117857600, 
    1117861200, 1117864800, 1117868400, 1117872000, 1117875600, 1117879200, 
    1117882800, 1117886400, 1117890000, 1117893600, 1117897200, 1117900800, 
    1117904400, 1117908000, 1117911600, 1117915200, 1117918800, 1117922400, 
    1117926000, 1117929600, 1117933200, 1117936800, 1117940400, 1117944000, 
    1117947600, 1117951200, 1117954800, 1117958400, 1117962000, 1117965600, 
    1117969200, 1117972800, 1117976400, 1117980000, 1117983600, 1117987200, 
    1117990800, 1117994400, 1117998000, 1118001600, 1118005200, 1118008800, 
    1118012400, 1118016000, 1118019600, 1118023200, 1118026800, 1118030400, 
    1118034000, 1118037600, 1118041200, 1118044800, 1118048400, 1118052000, 
    1118055600, 1118059200, 1118062800, 1118066400, 1118070000, 1118073600, 
    1118077200, 1118080800, 1118084400, 1118088000, 1118091600, 1118095200, 
    1118098800, 1118102400, 1118106000, 1118109600, 1118113200, 1118116800, 
    1118120400, 1118124000, 1118127600, 1118131200, 1118134800, 1118138400, 
    1118142000, 1118145600, 1118149200, 1118152800, 1118156400, 1118160000, 
    1118163600, 1118167200, 1118170800, 1118174400, 1118178000, 1118181600, 
    1118185200, 1118188800, 1118192400, 1118196000, 1118199600, 1118203200, 
    1118206800, 1118210400, 1118214000, 1118217600, 1118221200, 1118224800, 
    1118228400, 1118232000, 1118235600, 1118239200, 1118242800, 1118246400, 
    1118250000, 1118253600, 1118257200, 1118260800, 1118264400, 1118268000, 
    1118271600, 1118275200, 1118278800, 1118282400, 1118286000, 1118289600, 
    1118293200, 1118296800, 1118300400, 1118304000, 1118307600, 1118311200, 
    1118314800, 1118318400, 1118322000, 1118325600, 1118329200, 1118332800, 
    1118336400, 1118340000, 1118343600, 1118347200, 1118350800, 1118354400, 
    1118358000, 1118361600, 1118365200, 1118368800, 1118372400, 1118376000, 
    1118379600, 1118383200, 1118386800, 1118390400, 1118394000, 1118397600, 
    1118401200, 1118404800, 1118408400, 1118412000, 1118415600, 1118419200, 
    1118422800, 1118426400, 1118430000, 1118433600, 1118437200, 1118440800, 
    1118444400, 1118448000, 1118451600, 1118455200, 1118458800, 1118462400, 
    1118466000, 1118469600, 1118473200, 1118476800, 1118480400, 1118484000, 
    1118487600, 1118491200, 1118494800, 1118498400, 1118502000, 1118505600, 
    1118509200, 1118512800, 1118516400, 1118520000, 1118523600, 1118527200, 
    1118530800, 1118534400, 1118538000, 1118541600, 1118545200, 1118548800, 
    1118552400, 1118556000, 1118559600, 1118563200, 1118566800, 1118570400, 
    1118574000, 1118577600, 1118581200, 1118584800, 1118588400, 1118592000, 
    1118595600, 1118599200, 1118602800, 1118606400, 1118610000, 1118613600, 
    1118617200, 1118620800, 1118624400, 1118628000, 1118631600, 1118635200, 
    1118638800, 1118642400, 1118646000, 1118649600, 1118653200, 1118656800, 
    1118660400, 1118664000, 1118667600, 1118671200, 1118674800, 1118678400, 
    1118682000, 1118685600, 1118689200, 1118692800, 1118696400, 1118700000, 
    1118703600, 1118707200, 1118710800, 1118714400, 1118718000, 1118721600, 
    1118725200, 1118728800, 1118732400, 1118736000, 1118739600, 1118743200, 
    1118746800, 1118750400, 1118754000, 1118757600, 1118761200, 1118764800, 
    1118768400, 1118772000, 1118775600, 1118779200, 1118782800, 1118786400, 
    1118790000, 1118793600, 1118797200, 1118800800, 1118804400, 1118808000, 
    1118811600, 1118815200, 1118818800, 1118822400, 1118826000, 1118829600, 
    1118833200, 1118836800, 1118840400, 1118844000, 1118847600, 1118851200, 
    1118854800, 1118858400, 1118862000, 1118865600, 1118869200, 1118872800, 
    1118876400, 1118880000, 1118883600, 1118887200, 1118890800, 1118894400, 
    1118898000, 1118901600, 1118905200, 1118908800, 1118912400, 1118916000, 
    1118919600, 1118923200, 1118926800, 1118930400, 1118934000, 1118937600, 
    1118941200, 1118944800, 1118948400, 1118952000, 1118955600, 1118959200, 
    1118962800, 1118966400, 1118970000, 1118973600, 1118977200, 1118980800, 
    1118984400, 1118988000, 1118991600, 1118995200, 1118998800, 1119002400, 
    1119006000, 1119009600, 1119013200, 1119016800, 1119020400, 1119024000, 
    1119027600, 1119031200, 1119034800, 1119038400, 1119042000, 1119045600, 
    1119049200, 1119052800, 1119056400, 1119060000, 1119063600, 1119067200, 
    1119070800, 1119074400, 1119078000, 1119081600, 1119085200, 1119088800, 
    1119092400, 1119096000, 1119099600, 1119103200, 1119106800, 1119110400, 
    1119114000, 1119117600, 1119121200, 1119124800, 1119128400, 1119132000, 
    1119135600, 1119139200, 1119142800, 1119146400, 1119150000, 1119153600, 
    1119157200, 1119160800, 1119164400, 1119168000, 1119171600, 1119175200, 
    1119178800, 1119182400, 1119186000, 1119189600, 1119193200, 1119196800, 
    1119200400, 1119204000, 1119207600, 1119211200, 1119214800, 1119218400, 
    1119222000, 1119225600, 1119229200, 1119232800, 1119236400, 1119240000, 
    1119243600, 1119247200, 1119250800, 1119254400, 1119258000, 1119261600, 
    1119265200, 1119268800, 1119272400, 1119276000, 1119279600, 1119283200, 
    1119286800, 1119290400, 1119294000, 1119297600, 1119301200, 1119304800, 
    1119308400, 1119312000, 1119315600, 1119319200, 1119322800, 1119326400, 
    1119330000, 1119333600, 1119337200, 1119340800, 1119344400, 1119348000, 
    1119351600, 1119355200, 1119358800, 1119362400, 1119366000, 1119369600, 
    1119373200, 1119376800, 1119380400, 1119384000, 1119387600, 1119391200, 
    1119394800, 1119398400, 1119402000, 1119405600, 1119409200, 1119412800, 
    1119416400, 1119420000, 1119423600, 1119427200, 1119430800, 1119434400, 
    1119438000, 1119441600, 1119445200, 1119448800, 1119452400, 1119456000, 
    1119459600, 1119463200, 1119466800, 1119470400, 1119474000, 1119477600, 
    1119481200, 1119484800, 1119488400, 1119492000, 1119495600, 1119499200, 
    1119502800, 1119506400, 1119510000, 1119513600, 1119517200, 1119520800, 
    1119524400, 1119528000, 1119531600, 1119535200, 1119538800, 1119542400, 
    1119546000, 1119549600, 1119553200, 1119556800, 1119560400, 1119564000, 
    1119567600, 1119571200, 1119574800, 1119578400, 1119582000, 1119585600, 
    1119589200, 1119592800, 1119596400, 1119600000, 1119603600, 1119607200, 
    1119610800, 1119614400, 1119618000, 1119621600, 1119625200, 1119628800, 
    1119632400, 1119636000, 1119639600, 1119643200, 1119646800, 1119650400, 
    1119654000, 1119657600, 1119661200, 1119664800, 1119668400, 1119672000, 
    1119675600, 1119679200, 1119682800, 1119686400, 1119690000, 1119693600, 
    1119697200, 1119700800, 1119704400, 1119708000, 1119711600, 1119715200, 
    1119718800, 1119722400, 1119726000, 1119729600, 1119733200, 1119736800, 
    1119740400, 1119744000, 1119747600, 1119751200, 1119754800, 1119758400, 
    1119762000, 1119765600, 1119769200, 1119772800, 1119776400, 1119780000, 
    1119783600, 1119787200, 1119790800, 1119794400, 1119798000, 1119801600, 
    1119805200, 1119808800, 1119812400, 1119816000, 1119819600, 1119823200, 
    1119826800, 1119830400, 1119834000, 1119837600, 1119841200, 1119844800, 
    1119848400, 1119852000, 1119855600, 1119859200, 1119862800, 1119866400, 
    1119870000, 1119873600, 1119877200, 1119880800, 1119884400, 1119888000, 
    1119891600, 1119895200, 1119898800, 1119902400, 1119906000, 1119909600, 
    1119913200, 1119916800, 1119920400, 1119924000, 1119927600, 1119931200, 
    1119934800, 1119938400, 1119942000, 1119945600, 1119949200, 1119952800, 
    1119956400, 1119960000, 1119963600, 1119967200, 1119970800, 1119974400, 
    1119978000, 1119981600, 1119985200, 1119988800, 1119992400, 1119996000, 
    1119999600, 1120003200, 1120006800, 1120010400, 1120014000, 1120017600, 
    1120021200, 1120024800, 1120028400, 1120032000, 1120035600, 1120039200, 
    1120042800, 1120046400, 1120050000, 1120053600, 1120057200, 1120060800, 
    1120064400, 1120068000, 1120071600, 1120075200, 1120078800, 1120082400, 
    1120086000, 1120089600, 1120093200, 1120096800, 1120100400, 1120104000, 
    1120107600, 1120111200, 1120114800, 1120118400, 1120122000, 1120125600, 
    1120129200, 1120132800, 1120136400, 1120140000, 1120143600, 1120147200, 
    1120150800, 1120154400, 1120158000, 1120161600, 1120165200, 1120168800, 
    1120172400, 1120176000, 1120179600, 1120183200, 1120186800, 1120190400, 
    1120194000, 1120197600, 1120201200, 1120204800, 1120208400, 1120212000, 
    1120215600, 1120219200, 1120222800, 1120226400, 1120230000, 1120233600, 
    1120237200, 1120240800, 1120244400, 1120248000, 1120251600, 1120255200, 
    1120258800, 1120262400, 1120266000, 1120269600, 1120273200, 1120276800, 
    1120280400, 1120284000, 1120287600, 1120291200, 1120294800, 1120298400, 
    1120302000, 1120305600, 1120309200, 1120312800, 1120316400, 1120320000, 
    1120323600, 1120327200, 1120330800, 1120334400, 1120338000, 1120341600, 
    1120345200, 1120348800, 1120352400, 1120356000, 1120359600, 1120363200, 
    1120366800, 1120370400, 1120374000, 1120377600, 1120381200, 1120384800, 
    1120388400, 1120392000, 1120395600, 1120399200, 1120402800, 1120406400, 
    1120410000, 1120413600, 1120417200, 1120420800, 1120424400, 1120428000, 
    1120431600, 1120435200, 1120438800, 1120442400, 1120446000, 1120449600, 
    1120453200, 1120456800, 1120460400, 1120464000, 1120467600, 1120471200, 
    1120474800, 1120478400, 1120482000, 1120485600, 1120489200, 1120492800, 
    1120496400, 1120500000, 1120503600, 1120507200, 1120510800, 1120514400, 
    1120518000, 1120521600, 1120525200, 1120528800, 1120532400, 1120536000, 
    1120539600, 1120543200, 1120546800, 1120550400, 1120554000, 1120557600, 
    1120561200, 1120564800, 1120568400, 1120572000, 1120575600, 1120579200, 
    1120582800, 1120586400, 1120590000, 1120593600, 1120597200, 1120600800, 
    1120604400, 1120608000, 1120611600, 1120615200, 1120618800, 1120622400, 
    1120626000, 1120629600, 1120633200, 1120636800, 1120640400, 1120644000, 
    1120647600, 1120651200, 1120654800, 1120658400, 1120662000, 1120665600, 
    1120669200, 1120672800, 1120676400, 1120680000, 1120683600, 1120687200, 
    1120690800, 1120694400, 1120698000, 1120701600, 1120705200, 1120708800, 
    1120712400, 1120716000, 1120719600, 1120723200, 1120726800, 1120730400, 
    1120734000, 1120737600, 1120741200, 1120744800, 1120748400, 1120752000, 
    1120755600, 1120759200, 1120762800, 1120766400, 1120770000, 1120773600, 
    1120777200, 1120780800, 1120784400, 1120788000, 1120791600, 1120795200, 
    1120798800, 1120802400, 1120806000, 1120809600, 1120813200, 1120816800, 
    1120820400, 1120824000, 1120827600, 1120831200, 1120834800, 1120838400, 
    1120842000, 1120845600, 1120849200, 1120852800, 1120856400, 1120860000, 
    1120863600, 1120867200, 1120870800, 1120874400, 1120878000, 1120881600, 
    1120885200, 1120888800, 1120892400, 1120896000, 1120899600, 1120903200, 
    1120906800, 1120910400, 1120914000, 1120917600, 1120921200, 1120924800, 
    1120928400, 1120932000, 1120935600, 1120939200, 1120942800, 1120946400, 
    1120950000, 1120953600, 1120957200, 1120960800, 1120964400, 1120968000, 
    1120971600, 1120975200, 1120978800, 1120982400, 1120986000, 1120989600, 
    1120993200, 1120996800, 1121000400, 1121004000, 1121007600, 1121011200, 
    1121014800, 1121018400, 1121022000, 1121025600, 1121029200, 1121032800, 
    1121036400, 1121040000, 1121043600, 1121047200, 1121050800, 1121054400, 
    1121058000, 1121061600, 1121065200, 1121068800, 1121072400, 1121076000, 
    1121079600, 1121083200, 1121086800, 1121090400, 1121094000, 1121097600, 
    1121101200, 1121104800, 1121108400, 1121112000, 1121115600, 1121119200, 
    1121122800, 1121126400, 1121130000, 1121133600, 1121137200, 1121140800, 
    1121144400, 1121148000, 1121151600, 1121155200, 1121158800, 1121162400, 
    1121166000, 1121169600, 1121173200, 1121176800, 1121180400, 1121184000, 
    1121187600, 1121191200, 1121194800, 1121198400, 1121202000, 1121205600, 
    1121209200, 1121212800, 1121216400, 1121220000, 1121223600, 1121227200, 
    1121230800, 1121234400, 1121238000, 1121241600, 1121245200, 1121248800, 
    1121252400, 1121256000, 1121259600, 1121263200, 1121266800, 1121270400, 
    1121274000, 1121277600, 1121281200, 1121284800, 1121288400, 1121292000, 
    1121295600, 1121299200, 1121302800, 1121306400, 1121310000, 1121313600, 
    1121317200, 1121320800, 1121324400, 1121328000, 1121331600, 1121335200, 
    1121338800, 1121342400, 1121346000, 1121349600, 1121353200, 1121356800, 
    1121360400, 1121364000, 1121367600, 1121371200, 1121374800, 1121378400, 
    1121382000, 1121385600, 1121389200, 1121392800, 1121396400, 1121400000, 
    1121403600, 1121407200, 1121410800, 1121414400, 1121418000, 1121421600, 
    1121425200, 1121428800, 1121432400, 1121436000, 1121439600, 1121443200, 
    1121446800, 1121450400, 1121454000, 1121457600, 1121461200, 1121464800, 
    1121468400, 1121472000, 1121475600, 1121479200, 1121482800, 1121486400, 
    1121490000, 1121493600, 1121497200, 1121500800, 1121504400, 1121508000, 
    1121511600, 1121515200, 1121518800, 1121522400, 1121526000, 1121529600, 
    1121533200, 1121536800, 1121540400, 1121544000, 1121547600, 1121551200, 
    1121554800, 1121558400, 1121562000, 1121565600, 1121569200, 1121572800, 
    1121576400, 1121580000, 1121583600, 1121587200, 1121590800, 1121594400, 
    1121598000, 1121601600, 1121605200, 1121608800, 1121612400, 1121616000, 
    1121619600, 1121623200, 1121626800, 1121630400, 1121634000, 1121637600, 
    1121641200, 1121644800, 1121648400, 1121652000, 1121655600, 1121659200, 
    1121662800, 1121666400, 1121670000, 1121673600, 1121677200, 1121680800, 
    1121684400, 1121688000, 1121691600, 1121695200, 1121698800, 1121702400, 
    1121706000, 1121709600, 1121713200, 1121716800, 1121720400, 1121724000, 
    1121727600, 1121731200, 1121734800, 1121738400, 1121742000, 1121745600, 
    1121749200, 1121752800, 1121756400, 1121760000, 1121763600, 1121767200, 
    1121770800, 1121774400, 1121778000, 1121781600, 1121785200, 1121788800, 
    1121792400, 1121796000, 1121799600, 1121803200, 1121806800, 1121810400, 
    1121814000, 1121817600, 1121821200, 1121824800, 1121828400, 1121832000, 
    1121835600, 1121839200, 1121842800, 1121846400, 1121850000, 1121853600, 
    1121857200, 1121860800, 1121864400, 1121868000, 1121871600, 1121875200, 
    1121878800, 1121882400, 1121886000, 1121889600, 1121893200, 1121896800, 
    1121900400, 1121904000, 1121907600, 1121911200, 1121914800, 1121918400, 
    1121922000, 1121925600, 1121929200, 1121932800, 1121936400, 1121940000, 
    1121943600, 1121947200, 1121950800, 1121954400, 1121958000, 1121961600, 
    1121965200, 1121968800, 1121972400, 1121976000, 1121979600, 1121983200, 
    1121986800, 1121990400, 1121994000, 1121997600, 1122001200, 1122004800, 
    1122008400, 1122012000, 1122015600, 1122019200, 1122022800, 1122026400, 
    1122030000, 1122033600, 1122037200, 1122040800, 1122044400, 1122048000, 
    1122051600, 1122055200, 1122058800, 1122062400, 1122066000, 1122069600, 
    1122073200, 1122076800, 1122080400, 1122084000, 1122087600, 1122091200, 
    1122094800, 1122098400, 1122102000, 1122105600, 1122109200, 1122112800, 
    1122116400, 1122120000, 1122123600, 1122127200, 1122130800, 1122134400, 
    1122138000, 1122141600, 1122145200, 1122148800, 1122152400, 1122156000, 
    1122159600, 1122163200, 1122166800, 1122170400, 1122174000, 1122177600, 
    1122181200, 1122184800, 1122188400, 1122192000, 1122195600, 1122199200, 
    1122202800, 1122206400, 1122210000, 1122213600, 1122217200, 1122220800, 
    1122224400, 1122228000, 1122231600, 1122235200, 1122238800, 1122242400, 
    1122246000, 1122249600, 1122253200, 1122256800, 1122260400, 1122264000, 
    1122267600, 1122271200, 1122274800, 1122278400, 1122282000, 1122285600, 
    1122289200, 1122292800, 1122296400, 1122300000, 1122303600, 1122307200, 
    1122310800, 1122314400, 1122318000, 1122321600, 1122325200, 1122328800, 
    1122332400, 1122336000, 1122339600, 1122343200, 1122346800, 1122350400, 
    1122354000, 1122357600, 1122361200, 1122364800, 1122368400, 1122372000, 
    1122375600, 1122379200, 1122382800, 1122386400, 1122390000, 1122393600, 
    1122397200, 1122400800, 1122404400, 1122408000, 1122411600, 1122415200, 
    1122418800, 1122422400, 1122426000, 1122429600, 1122433200, 1122436800, 
    1122440400, 1122444000, 1122447600, 1122451200, 1122454800, 1122458400, 
    1122462000, 1122465600, 1122469200, 1122472800, 1122476400, 1122480000, 
    1122483600, 1122487200, 1122490800, 1122494400, 1122498000, 1122501600, 
    1122505200, 1122508800, 1122512400, 1122516000, 1122519600, 1122523200, 
    1122526800, 1122530400, 1122534000, 1122537600, 1122541200, 1122544800, 
    1122548400, 1122552000, 1122555600, 1122559200, 1122562800, 1122566400, 
    1122570000, 1122573600, 1122577200, 1122580800, 1122584400, 1122588000, 
    1122591600, 1122595200, 1122598800, 1122602400, 1122606000, 1122609600, 
    1122613200, 1122616800, 1122620400, 1122624000, 1122627600, 1122631200, 
    1122634800, 1122638400, 1122642000, 1122645600, 1122649200, 1122652800, 
    1122656400, 1122660000, 1122663600, 1122667200, 1122670800, 1122674400, 
    1122678000, 1122681600, 1122685200, 1122688800, 1122692400, 1122696000, 
    1122699600, 1122703200, 1122706800, 1122710400, 1122714000, 1122717600, 
    1122721200, 1122724800, 1122728400, 1122732000, 1122735600, 1122739200, 
    1122742800, 1122746400, 1122750000, 1122753600, 1122757200, 1122760800, 
    1122764400, 1122768000, 1122771600, 1122775200, 1122778800, 1122782400, 
    1122786000, 1122789600, 1122793200, 1122796800, 1122800400, 1122804000, 
    1122807600, 1122811200, 1122814800, 1122818400, 1122822000, 1122825600, 
    1122829200, 1122832800, 1122836400, 1122840000, 1122843600, 1122847200, 
    1122850800, 1122854400, 1122858000, 1122861600, 1122865200, 1122868800, 
    1122872400, 1122876000, 1122879600, 1122883200, 1122886800, 1122890400, 
    1122894000, 1122897600, 1122901200, 1122904800, 1122908400, 1122912000, 
    1122915600, 1122919200, 1122922800, 1122926400, 1122930000, 1122933600, 
    1122937200, 1122940800, 1122944400, 1122948000, 1122951600, 1122955200, 
    1122958800, 1122962400, 1122966000, 1122969600, 1122973200, 1122976800, 
    1122980400, 1122984000, 1122987600, 1122991200, 1122994800, 1122998400, 
    1123002000, 1123005600, 1123009200, 1123012800, 1123016400, 1123020000, 
    1123023600, 1123027200, 1123030800, 1123034400, 1123038000, 1123041600, 
    1123045200, 1123048800, 1123052400, 1123056000, 1123059600, 1123063200, 
    1123066800, 1123070400, 1123074000, 1123077600, 1123081200, 1123084800, 
    1123088400, 1123092000, 1123095600, 1123099200, 1123102800, 1123106400, 
    1123110000, 1123113600, 1123117200, 1123120800, 1123124400, 1123128000, 
    1123131600, 1123135200, 1123138800, 1123142400, 1123146000, 1123149600, 
    1123153200, 1123156800, 1123160400, 1123164000, 1123167600, 1123171200, 
    1123174800, 1123178400, 1123182000, 1123185600, 1123189200, 1123192800, 
    1123196400, 1123200000, 1123203600, 1123207200, 1123210800, 1123214400, 
    1123218000, 1123221600, 1123225200, 1123228800, 1123232400, 1123236000, 
    1123239600, 1123243200, 1123246800, 1123250400, 1123254000, 1123257600, 
    1123261200, 1123264800, 1123268400, 1123272000, 1123275600, 1123279200, 
    1123282800, 1123286400, 1123290000, 1123293600, 1123297200, 1123300800, 
    1123304400, 1123308000, 1123311600, 1123315200, 1123318800, 1123322400, 
    1123326000, 1123329600, 1123333200, 1123336800, 1123340400, 1123344000, 
    1123347600, 1123351200, 1123354800, 1123358400, 1123362000, 1123365600, 
    1123369200, 1123372800, 1123376400, 1123380000, 1123383600, 1123387200, 
    1123390800, 1123394400, 1123398000, 1123401600, 1123405200, 1123408800, 
    1123412400, 1123416000, 1123419600, 1123423200, 1123426800, 1123430400, 
    1123434000, 1123437600, 1123441200, 1123444800, 1123448400, 1123452000, 
    1123455600, 1123459200, 1123462800, 1123466400, 1123470000, 1123473600, 
    1123477200, 1123480800, 1123484400, 1123488000, 1123491600, 1123495200, 
    1123498800, 1123502400, 1123506000, 1123509600, 1123513200, 1123516800, 
    1123520400, 1123524000, 1123527600, 1123531200, 1123534800, 1123538400, 
    1123542000, 1123545600, 1123549200, 1123552800, 1123556400, 1123560000, 
    1123563600, 1123567200, 1123570800, 1123574400, 1123578000, 1123581600, 
    1123585200, 1123588800, 1123592400, 1123596000, 1123599600, 1123603200, 
    1123606800, 1123610400, 1123614000, 1123617600, 1123621200, 1123624800, 
    1123628400, 1123632000, 1123635600, 1123639200, 1123642800, 1123646400, 
    1123650000, 1123653600, 1123657200, 1123660800, 1123664400, 1123668000, 
    1123671600, 1123675200, 1123678800, 1123682400, 1123686000, 1123689600, 
    1123693200, 1123696800, 1123700400, 1123704000, 1123707600, 1123711200, 
    1123714800, 1123718400, 1123722000, 1123725600, 1123729200, 1123732800, 
    1123736400, 1123740000, 1123743600, 1123747200, 1123750800, 1123754400, 
    1123758000, 1123761600, 1123765200, 1123768800, 1123772400, 1123776000, 
    1123779600, 1123783200, 1123786800, 1123790400, 1123794000, 1123797600, 
    1123801200, 1123804800, 1123808400, 1123812000, 1123815600, 1123819200, 
    1123822800, 1123826400, 1123830000, 1123833600, 1123837200, 1123840800, 
    1123844400, 1123848000, 1123851600, 1123855200, 1123858800, 1123862400, 
    1123866000, 1123869600, 1123873200, 1123876800, 1123880400, 1123884000, 
    1123887600, 1123891200, 1123894800, 1123898400, 1123902000, 1123905600, 
    1123909200, 1123912800, 1123916400, 1123920000, 1123923600, 1123927200, 
    1123930800, 1123934400, 1123938000, 1123941600, 1123945200, 1123948800, 
    1123952400, 1123956000, 1123959600, 1123963200, 1123966800, 1123970400, 
    1123974000, 1123977600, 1123981200, 1123984800, 1123988400, 1123992000, 
    1123995600, 1123999200, 1124002800, 1124006400, 1124010000, 1124013600, 
    1124017200, 1124020800, 1124024400, 1124028000, 1124031600, 1124035200, 
    1124038800, 1124042400, 1124046000, 1124049600, 1124053200, 1124056800, 
    1124060400, 1124064000, 1124067600, 1124071200, 1124074800, 1124078400, 
    1124082000, 1124085600, 1124089200, 1124092800, 1124096400, 1124100000, 
    1124103600, 1124107200, 1124110800, 1124114400, 1124118000, 1124121600, 
    1124125200, 1124128800, 1124132400, 1124136000, 1124139600, 1124143200, 
    1124146800, 1124150400, 1124154000, 1124157600, 1124161200, 1124164800, 
    1124168400, 1124172000, 1124175600, 1124179200, 1124182800, 1124186400, 
    1124190000, 1124193600, 1124197200, 1124200800, 1124204400, 1124208000, 
    1124211600, 1124215200, 1124218800, 1124222400, 1124226000, 1124229600, 
    1124233200, 1124236800, 1124240400, 1124244000, 1124247600, 1124251200, 
    1124254800, 1124258400, 1124262000, 1124265600, 1124269200, 1124272800, 
    1124276400, 1124280000, 1124283600, 1124287200, 1124290800, 1124294400, 
    1124298000, 1124301600, 1124305200, 1124308800, 1124312400, 1124316000, 
    1124319600, 1124323200, 1124326800, 1124330400, 1124334000, 1124337600, 
    1124341200, 1124344800, 1124348400, 1124352000, 1124355600, 1124359200, 
    1124362800, 1124366400, 1124370000, 1124373600, 1124377200, 1124380800, 
    1124384400, 1124388000, 1124391600, 1124395200, 1124398800, 1124402400, 
    1124406000, 1124409600, 1124413200, 1124416800, 1124420400, 1124424000, 
    1124427600, 1124431200, 1124434800, 1124438400, 1124442000, 1124445600, 
    1124449200, 1124452800, 1124456400, 1124460000, 1124463600, 1124467200, 
    1124470800, 1124474400, 1124478000, 1124481600, 1124485200, 1124488800, 
    1124492400, 1124496000, 1124499600, 1124503200, 1124506800, 1124510400, 
    1124514000, 1124517600, 1124521200, 1124524800, 1124528400, 1124532000, 
    1124535600, 1124539200, 1124542800, 1124546400, 1124550000, 1124553600, 
    1124557200, 1124560800, 1124564400, 1124568000, 1124571600, 1124575200, 
    1124578800, 1124582400, 1124586000, 1124589600, 1124593200, 1124596800, 
    1124600400, 1124604000, 1124607600, 1124611200, 1124614800, 1124618400, 
    1124622000, 1124625600, 1124629200, 1124632800, 1124636400, 1124640000, 
    1124643600, 1124647200, 1124650800, 1124654400, 1124658000, 1124661600, 
    1124665200, 1124668800, 1124672400, 1124676000, 1124679600, 1124683200, 
    1124686800, 1124690400, 1124694000, 1124697600, 1124701200, 1124704800, 
    1124708400, 1124712000, 1124715600, 1124719200, 1124722800, 1124726400, 
    1124730000, 1124733600, 1124737200, 1124740800, 1124744400, 1124748000, 
    1124751600, 1124755200, 1124758800, 1124762400, 1124766000, 1124769600, 
    1124773200, 1124776800, 1124780400, 1124784000, 1124787600, 1124791200, 
    1124794800, 1124798400, 1124802000, 1124805600, 1124809200, 1124812800, 
    1124816400, 1124820000, 1124823600, 1124827200, 1124830800, 1124834400, 
    1124838000, 1124841600, 1124845200, 1124848800, 1124852400, 1124856000, 
    1124859600, 1124863200, 1124866800, 1124870400, 1124874000, 1124877600, 
    1124881200, 1124884800, 1124888400, 1124892000, 1124895600, 1124899200, 
    1124902800, 1124906400, 1124910000, 1124913600, 1124917200, 1124920800, 
    1124924400, 1124928000, 1124931600, 1124935200, 1124938800, 1124942400, 
    1124946000, 1124949600, 1124953200, 1124956800, 1124960400, 1124964000, 
    1124967600, 1124971200, 1124974800, 1124978400, 1124982000, 1124985600, 
    1124989200, 1124992800, 1124996400, 1125000000, 1125003600, 1125007200, 
    1125010800, 1125014400, 1125018000, 1125021600, 1125025200, 1125028800, 
    1125032400, 1125036000, 1125039600, 1125043200, 1125046800, 1125050400, 
    1125054000, 1125057600, 1125061200, 1125064800, 1125068400, 1125072000, 
    1125075600, 1125079200, 1125082800, 1125086400, 1125090000, 1125093600, 
    1125097200, 1125100800, 1125104400, 1125108000, 1125111600, 1125115200, 
    1125118800, 1125122400, 1125126000, 1125129600, 1125133200, 1125136800, 
    1125140400, 1125144000, 1125147600, 1125151200, 1125154800, 1125158400, 
    1125162000, 1125165600, 1125169200, 1125172800, 1125176400, 1125180000, 
    1125183600, 1125187200, 1125190800, 1125194400, 1125198000, 1125201600, 
    1125205200, 1125208800, 1125212400, 1125216000, 1125219600, 1125223200, 
    1125226800, 1125230400, 1125234000, 1125237600, 1125241200, 1125244800, 
    1125248400, 1125252000, 1125255600, 1125259200, 1125262800, 1125266400, 
    1125270000, 1125273600, 1125277200, 1125280800, 1125284400, 1125288000, 
    1125291600, 1125295200, 1125298800, 1125302400, 1125306000, 1125309600, 
    1125313200, 1125316800, 1125320400, 1125324000, 1125327600, 1125331200, 
    1125334800, 1125338400, 1125342000, 1125345600, 1125349200, 1125352800, 
    1125356400, 1125360000, 1125363600, 1125367200, 1125370800, 1125374400, 
    1125378000, 1125381600, 1125385200, 1125388800, 1125392400, 1125396000, 
    1125399600, 1125403200, 1125406800, 1125410400, 1125414000, 1125417600, 
    1125421200, 1125424800, 1125428400, 1125432000, 1125435600, 1125439200, 
    1125442800, 1125446400, 1125450000, 1125453600, 1125457200, 1125460800, 
    1125464400, 1125468000, 1125471600, 1125475200, 1125478800, 1125482400, 
    1125486000, 1125489600, 1125493200, 1125496800, 1125500400, 1125504000, 
    1125507600, 1125511200, 1125514800, 1125518400, 1125522000, 1125525600, 
    1125529200, 1125532800, 1125536400, 1125540000, 1125543600, 1125547200, 
    1125550800, 1125554400, 1125558000, 1125561600, 1125565200, 1125568800, 
    1125572400, 1125576000, 1125579600, 1125583200, 1125586800, 1125590400, 
    1125594000, 1125597600, 1125601200, 1125604800, 1125608400, 1125612000, 
    1125615600, 1125619200, 1125622800, 1125626400, 1125630000, 1125633600, 
    1125637200, 1125640800, 1125644400, 1125648000, 1125651600, 1125655200, 
    1125658800, 1125662400, 1125666000, 1125669600, 1125673200, 1125676800, 
    1125680400, 1125684000, 1125687600, 1125691200, 1125694800, 1125698400, 
    1125702000, 1125705600, 1125709200, 1125712800, 1125716400, 1125720000, 
    1125723600, 1125727200, 1125730800, 1125734400, 1125738000, 1125741600, 
    1125745200, 1125748800, 1125752400, 1125756000, 1125759600, 1125763200, 
    1125766800, 1125770400, 1125774000, 1125777600, 1125781200, 1125784800, 
    1125788400, 1125792000, 1125795600, 1125799200, 1125802800, 1125806400, 
    1125810000, 1125813600, 1125817200, 1125820800, 1125824400, 1125828000, 
    1125831600, 1125835200, 1125838800, 1125842400, 1125846000, 1125849600, 
    1125853200, 1125856800, 1125860400, 1125864000, 1125867600, 1125871200, 
    1125874800, 1125878400, 1125882000, 1125885600, 1125889200, 1125892800, 
    1125896400, 1125900000, 1125903600, 1125907200, 1125910800, 1125914400, 
    1125918000, 1125921600, 1125925200, 1125928800, 1125932400, 1125936000, 
    1125939600, 1125943200, 1125946800, 1125950400, 1125954000, 1125957600, 
    1125961200, 1125964800, 1125968400, 1125972000, 1125975600, 1125979200, 
    1125982800, 1125986400, 1125990000, 1125993600, 1125997200, 1126000800, 
    1126004400, 1126008000, 1126011600, 1126015200, 1126018800, 1126022400, 
    1126026000, 1126029600, 1126033200, 1126036800, 1126040400, 1126044000, 
    1126047600, 1126051200, 1126054800, 1126058400, 1126062000, 1126065600, 
    1126069200, 1126072800, 1126076400, 1126080000, 1126083600, 1126087200, 
    1126090800, 1126094400, 1126098000, 1126101600, 1126105200, 1126108800, 
    1126112400, 1126116000, 1126119600, 1126123200, 1126126800, 1126130400, 
    1126134000, 1126137600, 1126141200, 1126144800, 1126148400, 1126152000, 
    1126155600, 1126159200, 1126162800, 1126166400, 1126170000, 1126173600, 
    1126177200, 1126180800, 1126184400, 1126188000, 1126191600, 1126195200, 
    1126198800, 1126202400, 1126206000, 1126209600, 1126213200, 1126216800, 
    1126220400, 1126224000, 1126227600, 1126231200, 1126234800, 1126238400, 
    1126242000, 1126245600, 1126249200, 1126252800, 1126256400, 1126260000, 
    1126263600, 1126267200, 1126270800, 1126274400, 1126278000, 1126281600, 
    1126285200, 1126288800, 1126292400, 1126296000, 1126299600, 1126303200, 
    1126306800, 1126310400, 1126314000, 1126317600, 1126321200, 1126324800, 
    1126328400, 1126332000, 1126335600, 1126339200, 1126342800, 1126346400, 
    1126350000, 1126353600, 1126357200, 1126360800, 1126364400, 1126368000, 
    1126371600, 1126375200, 1126378800, 1126382400, 1126386000, 1126389600, 
    1126393200, 1126396800, 1126400400, 1126404000, 1126407600, 1126411200, 
    1126414800, 1126418400, 1126422000, 1126425600, 1126429200, 1126432800, 
    1126436400, 1126440000, 1126443600, 1126447200, 1126450800, 1126454400, 
    1126458000, 1126461600, 1126465200, 1126468800, 1126472400, 1126476000, 
    1126479600, 1126483200, 1126486800, 1126490400, 1126494000, 1126497600, 
    1126501200, 1126504800, 1126508400, 1126512000, 1126515600, 1126519200, 
    1126522800, 1126526400, 1126530000, 1126533600, 1126537200, 1126540800, 
    1126544400, 1126548000, 1126551600, 1126555200, 1126558800, 1126562400, 
    1126566000, 1126569600, 1126573200, 1126576800, 1126580400, 1126584000, 
    1126587600, 1126591200, 1126594800, 1126598400, 1126602000, 1126605600, 
    1126609200, 1126612800, 1126616400, 1126620000, 1126623600, 1126627200, 
    1126630800, 1126634400, 1126638000, 1126641600, 1126645200, 1126648800, 
    1126652400, 1126656000, 1126659600, 1126663200, 1126666800, 1126670400, 
    1126674000, 1126677600, 1126681200, 1126684800, 1126688400, 1126692000, 
    1126695600, 1126699200, 1126702800, 1126706400, 1126710000, 1126713600, 
    1126717200, 1126720800, 1126724400, 1126728000, 1126731600, 1126735200, 
    1126738800, 1126742400, 1126746000, 1126749600, 1126753200, 1126756800, 
    1126760400, 1126764000, 1126767600, 1126771200, 1126774800, 1126778400, 
    1126782000, 1126785600, 1126789200, 1126792800, 1126796400, 1126800000, 
    1126803600, 1126807200, 1126810800, 1126814400, 1126818000, 1126821600, 
    1126825200, 1126828800, 1126832400, 1126836000, 1126839600, 1126843200, 
    1126846800, 1126850400, 1126854000, 1126857600, 1126861200, 1126864800, 
    1126868400, 1126872000, 1126875600, 1126879200, 1126882800, 1126886400, 
    1126890000, 1126893600, 1126897200, 1126900800, 1126904400, 1126908000, 
    1126911600, 1126915200, 1126918800, 1126922400, 1126926000, 1126929600, 
    1126933200, 1126936800, 1126940400, 1126944000, 1126947600, 1126951200, 
    1126954800, 1126958400, 1126962000, 1126965600, 1126969200, 1126972800, 
    1126976400, 1126980000, 1126983600, 1126987200, 1126990800, 1126994400, 
    1126998000, 1127001600, 1127005200, 1127008800, 1127012400, 1127016000, 
    1127019600, 1127023200, 1127026800, 1127030400, 1127034000, 1127037600, 
    1127041200, 1127044800, 1127048400, 1127052000, 1127055600, 1127059200, 
    1127062800, 1127066400, 1127070000, 1127073600, 1127077200, 1127080800, 
    1127084400, 1127088000, 1127091600, 1127095200, 1127098800, 1127102400, 
    1127106000, 1127109600, 1127113200, 1127116800, 1127120400, 1127124000, 
    1127127600, 1127131200, 1127134800, 1127138400, 1127142000, 1127145600, 
    1127149200, 1127152800, 1127156400, 1127160000, 1127163600, 1127167200, 
    1127170800, 1127174400, 1127178000, 1127181600, 1127185200, 1127188800, 
    1127192400, 1127196000, 1127199600, 1127203200, 1127206800, 1127210400, 
    1127214000, 1127217600, 1127221200, 1127224800, 1127228400, 1127232000, 
    1127235600, 1127239200, 1127242800, 1127246400, 1127250000, 1127253600, 
    1127257200, 1127260800, 1127264400, 1127268000, 1127271600, 1127275200, 
    1127278800, 1127282400, 1127286000, 1127289600, 1127293200, 1127296800, 
    1127300400, 1127304000, 1127307600, 1127311200, 1127314800, 1127318400, 
    1127322000, 1127325600, 1127329200, 1127332800, 1127336400, 1127340000, 
    1127343600, 1127347200, 1127350800, 1127354400, 1127358000, 1127361600, 
    1127365200, 1127368800, 1127372400, 1127376000, 1127379600, 1127383200, 
    1127386800, 1127390400, 1127394000, 1127397600, 1127401200, 1127404800, 
    1127408400, 1127412000, 1127415600, 1127419200, 1127422800, 1127426400, 
    1127430000, 1127433600, 1127437200, 1127440800, 1127444400, 1127448000, 
    1127451600, 1127455200, 1127458800, 1127462400, 1127466000, 1127469600, 
    1127473200, 1127476800, 1127480400, 1127484000, 1127487600, 1127491200, 
    1127494800, 1127498400, 1127502000, 1127505600, 1127509200, 1127512800, 
    1127516400, 1127520000, 1127523600, 1127527200, 1127530800, 1127534400, 
    1127538000, 1127541600, 1127545200, 1127548800, 1127552400, 1127556000, 
    1127559600, 1127563200, 1127566800, 1127570400, 1127574000, 1127577600, 
    1127581200, 1127584800, 1127588400, 1127592000, 1127595600, 1127599200, 
    1127602800, 1127606400, 1127610000, 1127613600, 1127617200, 1127620800, 
    1127624400, 1127628000, 1127631600, 1127635200, 1127638800, 1127642400, 
    1127646000, 1127649600, 1127653200, 1127656800, 1127660400, 1127664000, 
    1127667600, 1127671200, 1127674800, 1127678400, 1127682000, 1127685600, 
    1127689200, 1127692800, 1127696400, 1127700000, 1127703600, 1127707200, 
    1127710800, 1127714400, 1127718000, 1127721600, 1127725200, 1127728800, 
    1127732400, 1127736000, 1127739600, 1127743200, 1127746800, 1127750400, 
    1127754000, 1127757600, 1127761200, 1127764800, 1127768400, 1127772000, 
    1127775600, 1127779200, 1127782800, 1127786400, 1127790000, 1127793600, 
    1127797200, 1127800800, 1127804400, 1127808000, 1127811600, 1127815200, 
    1127818800, 1127822400, 1127826000, 1127829600, 1127833200, 1127836800, 
    1127840400, 1127844000, 1127847600, 1127851200, 1127854800, 1127858400, 
    1127862000, 1127865600, 1127869200, 1127872800, 1127876400, 1127880000, 
    1127883600, 1127887200, 1127890800, 1127894400, 1127898000, 1127901600, 
    1127905200, 1127908800, 1127912400, 1127916000, 1127919600, 1127923200, 
    1127926800, 1127930400, 1127934000, 1127937600, 1127941200, 1127944800, 
    1127948400, 1127952000, 1127955600, 1127959200, 1127962800, 1127966400, 
    1127970000, 1127973600, 1127977200, 1127980800, 1127984400, 1127988000, 
    1127991600, 1127995200, 1127998800, 1128002400, 1128006000, 1128009600, 
    1128013200, 1128016800, 1128020400, 1128024000, 1128027600, 1128031200, 
    1128034800, 1128038400, 1128042000, 1128045600, 1128049200, 1128052800, 
    1128056400, 1128060000, 1128063600, 1128067200, 1128070800, 1128074400, 
    1128078000, 1128081600, 1128085200, 1128088800, 1128092400, 1128096000, 
    1128099600, 1128103200, 1128106800, 1128110400, 1128114000, 1128117600, 
    1128121200, 1128124800, 1128128400, 1128132000, 1128135600, 1128139200, 
    1128142800, 1128146400, 1128150000, 1128153600, 1128157200, 1128160800, 
    1128164400, 1128168000, 1128171600, 1128175200, 1128178800, 1128182400, 
    1128186000, 1128189600, 1128193200, 1128196800, 1128200400, 1128204000, 
    1128207600, 1128211200, 1128214800, 1128218400, 1128222000, 1128225600, 
    1128229200, 1128232800, 1128236400, 1128240000, 1128243600, 1128247200, 
    1128250800, 1128254400, 1128258000, 1128261600, 1128265200, 1128268800, 
    1128272400, 1128276000, 1128279600, 1128283200, 1128286800, 1128290400, 
    1128294000, 1128297600, 1128301200, 1128304800, 1128308400, 1128312000, 
    1128315600, 1128319200, 1128322800, 1128326400, 1128330000, 1128333600, 
    1128337200, 1128340800, 1128344400, 1128348000, 1128351600, 1128355200, 
    1128358800, 1128362400, 1128366000, 1128369600, 1128373200, 1128376800, 
    1128380400, 1128384000, 1128387600, 1128391200, 1128394800, 1128398400, 
    1128402000, 1128405600, 1128409200, 1128412800, 1128416400, 1128420000, 
    1128423600, 1128427200, 1128430800, 1128434400, 1128438000, 1128441600, 
    1128445200, 1128448800, 1128452400, 1128456000, 1128459600, 1128463200, 
    1128466800, 1128470400, 1128474000, 1128477600, 1128481200, 1128484800, 
    1128488400, 1128492000, 1128495600, 1128499200, 1128502800, 1128506400, 
    1128510000, 1128513600, 1128517200, 1128520800, 1128524400, 1128528000, 
    1128531600, 1128535200, 1128538800, 1128542400, 1128546000, 1128549600, 
    1128553200, 1128556800, 1128560400, 1128564000, 1128567600, 1128571200, 
    1128574800, 1128578400, 1128582000, 1128585600, 1128589200, 1128592800, 
    1128596400, 1128600000, 1128603600, 1128607200, 1128610800, 1128614400, 
    1128618000, 1128621600, 1128625200, 1128628800, 1128632400, 1128636000, 
    1128639600, 1128643200, 1128646800, 1128650400, 1128654000, 1128657600, 
    1128661200, 1128664800, 1128668400, 1128672000, 1128675600, 1128679200, 
    1128682800, 1128686400, 1128690000, 1128693600, 1128697200, 1128700800, 
    1128704400, 1128708000, 1128711600, 1128715200, 1128718800, 1128722400, 
    1128726000, 1128729600, 1128733200, 1128736800, 1128740400, 1128744000, 
    1128747600, 1128751200, 1128754800, 1128758400, 1128762000, 1128765600, 
    1128769200, 1128772800, 1128776400, 1128780000, 1128783600, 1128787200, 
    1128790800, 1128794400, 1128798000, 1128801600, 1128805200, 1128808800, 
    1128812400, 1128816000, 1128819600, 1128823200, 1128826800, 1128830400, 
    1128834000, 1128837600, 1128841200, 1128844800, 1128848400, 1128852000, 
    1128855600, 1128859200, 1128862800, 1128866400, 1128870000, 1128873600, 
    1128877200, 1128880800, 1128884400, 1128888000, 1128891600, 1128895200, 
    1128898800, 1128902400, 1128906000, 1128909600, 1128913200, 1128916800, 
    1128920400, 1128924000, 1128927600, 1128931200, 1128934800, 1128938400, 
    1128942000, 1128945600, 1128949200, 1128952800, 1128956400, 1128960000, 
    1128963600, 1128967200, 1128970800, 1128974400, 1128978000, 1128981600, 
    1128985200, 1128988800, 1128992400, 1128996000, 1128999600, 1129003200, 
    1129006800, 1129010400, 1129014000, 1129017600, 1129021200, 1129024800, 
    1129028400, 1129032000, 1129035600, 1129039200, 1129042800, 1129046400, 
    1129050000, 1129053600, 1129057200, 1129060800, 1129064400, 1129068000, 
    1129071600, 1129075200, 1129078800, 1129082400, 1129086000, 1129089600, 
    1129093200, 1129096800, 1129100400, 1129104000, 1129107600, 1129111200, 
    1129114800, 1129118400, 1129122000, 1129125600, 1129129200, 1129132800, 
    1129136400, 1129140000, 1129143600, 1129147200, 1129150800, 1129154400, 
    1129158000, 1129161600, 1129165200, 1129168800, 1129172400, 1129176000, 
    1129179600, 1129183200, 1129186800, 1129190400, 1129194000, 1129197600, 
    1129201200, 1129204800, 1129208400, 1129212000, 1129215600, 1129219200, 
    1129222800, 1129226400, 1129230000, 1129233600, 1129237200, 1129240800, 
    1129244400, 1129248000, 1129251600, 1129255200, 1129258800, 1129262400, 
    1129266000, 1129269600, 1129273200, 1129276800, 1129280400, 1129284000, 
    1129287600, 1129291200, 1129294800, 1129298400, 1129302000, 1129305600, 
    1129309200, 1129312800, 1129316400, 1129320000, 1129323600, 1129327200, 
    1129330800, 1129334400, 1129338000, 1129341600, 1129345200, 1129348800, 
    1129352400, 1129356000, 1129359600, 1129363200, 1129366800, 1129370400, 
    1129374000, 1129377600, 1129381200, 1129384800, 1129388400, 1129392000, 
    1129395600, 1129399200, 1129402800, 1129406400, 1129410000, 1129413600, 
    1129417200, 1129420800, 1129424400, 1129428000, 1129431600, 1129435200, 
    1129438800, 1129442400, 1129446000, 1129449600, 1129453200, 1129456800, 
    1129460400, 1129464000, 1129467600, 1129471200, 1129474800, 1129478400, 
    1129482000, 1129485600, 1129489200, 1129492800, 1129496400, 1129500000, 
    1129503600, 1129507200, 1129510800, 1129514400, 1129518000, 1129521600, 
    1129525200, 1129528800, 1129532400, 1129536000, 1129539600, 1129543200, 
    1129546800, 1129550400, 1129554000, 1129557600, 1129561200, 1129564800, 
    1129568400, 1129572000, 1129575600, 1129579200, 1129582800, 1129586400, 
    1129590000, 1129593600, 1129597200, 1129600800, 1129604400, 1129608000, 
    1129611600, 1129615200, 1129618800, 1129622400, 1129626000, 1129629600, 
    1129633200, 1129636800, 1129640400, 1129644000, 1129647600, 1129651200, 
    1129654800, 1129658400, 1129662000, 1129665600, 1129669200, 1129672800, 
    1129676400, 1129680000, 1129683600, 1129687200, 1129690800, 1129694400, 
    1129698000, 1129701600, 1129705200, 1129708800, 1129712400, 1129716000, 
    1129719600, 1129723200, 1129726800, 1129730400, 1129734000, 1129737600, 
    1129741200, 1129744800, 1129748400, 1129752000, 1129755600, 1129759200, 
    1129762800, 1129766400, 1129770000, 1129773600, 1129777200, 1129780800, 
    1129784400, 1129788000, 1129791600, 1129795200, 1129798800, 1129802400, 
    1129806000, 1129809600, 1129813200, 1129816800, 1129820400, 1129824000, 
    1129827600, 1129831200, 1129834800, 1129838400, 1129842000, 1129845600, 
    1129849200, 1129852800, 1129856400, 1129860000, 1129863600, 1129867200, 
    1129870800, 1129874400, 1129878000, 1129881600, 1129885200, 1129888800, 
    1129892400, 1129896000, 1129899600, 1129903200, 1129906800, 1129910400, 
    1129914000, 1129917600, 1129921200, 1129924800, 1129928400, 1129932000, 
    1129935600, 1129939200, 1129942800, 1129946400, 1129950000, 1129953600, 
    1129957200, 1129960800, 1129964400, 1129968000, 1129971600, 1129975200, 
    1129978800, 1129982400, 1129986000, 1129989600, 1129993200, 1129996800, 
    1130000400, 1130004000, 1130007600, 1130011200, 1130014800, 1130018400, 
    1130022000, 1130025600, 1130029200, 1130032800, 1130036400, 1130040000, 
    1130043600, 1130047200, 1130050800, 1130054400, 1130058000, 1130061600, 
    1130065200, 1130068800, 1130072400, 1130076000, 1130079600, 1130083200, 
    1130086800, 1130090400, 1130094000, 1130097600, 1130101200, 1130104800, 
    1130108400, 1130112000, 1130115600, 1130119200, 1130122800, 1130126400, 
    1130130000, 1130133600, 1130137200, 1130140800, 1130144400, 1130148000, 
    1130151600, 1130155200, 1130158800, 1130162400, 1130166000, 1130169600, 
    1130173200, 1130176800, 1130180400, 1130184000, 1130187600, 1130191200, 
    1130194800, 1130198400, 1130202000, 1130205600, 1130209200, 1130212800, 
    1130216400, 1130220000, 1130223600, 1130227200, 1130230800, 1130234400, 
    1130238000, 1130241600, 1130245200, 1130248800, 1130252400, 1130256000, 
    1130259600, 1130263200, 1130266800, 1130270400, 1130274000, 1130277600, 
    1130281200, 1130284800, 1130288400, 1130292000, 1130295600, 1130299200, 
    1130302800, 1130306400, 1130310000, 1130313600, 1130317200, 1130320800, 
    1130324400, 1130328000, 1130331600, 1130335200, 1130338800, 1130342400, 
    1130346000, 1130349600, 1130353200, 1130356800, 1130360400, 1130364000, 
    1130367600, 1130371200, 1130374800, 1130378400, 1130382000, 1130385600, 
    1130389200, 1130392800, 1130396400, 1130400000, 1130403600, 1130407200, 
    1130410800, 1130414400, 1130418000, 1130421600, 1130425200, 1130428800, 
    1130432400, 1130436000, 1130439600, 1130443200, 1130446800, 1130450400, 
    1130454000, 1130457600, 1130461200, 1130464800, 1130468400, 1130472000, 
    1130475600, 1130479200, 1130482800, 1130486400, 1130490000, 1130493600, 
    1130497200, 1130500800, 1130504400, 1130508000, 1130511600, 1130515200, 
    1130518800, 1130522400, 1130526000, 1130529600, 1130533200, 1130536800, 
    1130540400, 1130544000, 1130547600, 1130551200, 1130554800, 1130558400, 
    1130562000, 1130565600, 1130569200, 1130572800, 1130576400, 1130580000, 
    1130583600, 1130587200, 1130590800, 1130594400, 1130598000, 1130601600, 
    1130605200, 1130608800, 1130612400, 1130616000, 1130619600, 1130623200, 
    1130626800, 1130630400, 1130634000, 1130637600, 1130641200, 1130644800, 
    1130648400, 1130652000, 1130655600, 1130659200, 1130662800, 1130666400, 
    1130670000, 1130673600, 1130677200, 1130680800, 1130684400, 1130688000, 
    1130691600, 1130695200, 1130698800, 1130702400, 1130706000, 1130709600, 
    1130713200, 1130716800, 1130720400, 1130724000, 1130727600, 1130731200, 
    1130734800, 1130738400, 1130742000, 1130745600, 1130749200, 1130752800, 
    1130756400, 1130760000, 1130763600, 1130767200, 1130770800, 1130774400, 
    1130778000, 1130781600, 1130785200, 1130788800, 1130792400, 1130796000, 
    1130799600, 1130803200, 1130806800, 1130810400, 1130814000, 1130817600, 
    1130821200, 1130824800, 1130828400, 1130832000, 1130835600, 1130839200, 
    1130842800, 1130846400, 1130850000, 1130853600, 1130857200, 1130860800, 
    1130864400, 1130868000, 1130871600, 1130875200, 1130878800, 1130882400, 
    1130886000, 1130889600, 1130893200, 1130896800, 1130900400, 1130904000, 
    1130907600, 1130911200, 1130914800, 1130918400, 1130922000, 1130925600, 
    1130929200, 1130932800, 1130936400, 1130940000, 1130943600, 1130947200, 
    1130950800, 1130954400, 1130958000, 1130961600, 1130965200, 1130968800, 
    1130972400, 1130976000, 1130979600, 1130983200, 1130986800, 1130990400, 
    1130994000, 1130997600, 1131001200, 1131004800, 1131008400, 1131012000, 
    1131015600, 1131019200, 1131022800, 1131026400, 1131030000, 1131033600, 
    1131037200, 1131040800, 1131044400, 1131048000, 1131051600, 1131055200, 
    1131058800, 1131062400, 1131066000, 1131069600, 1131073200, 1131076800, 
    1131080400, 1131084000, 1131087600, 1131091200, 1131094800, 1131098400, 
    1131102000, 1131105600, 1131109200, 1131112800, 1131116400, 1131120000, 
    1131123600, 1131127200, 1131130800, 1131134400, 1131138000, 1131141600, 
    1131145200, 1131148800, 1131152400, 1131156000, 1131159600, 1131163200, 
    1131166800, 1131170400, 1131174000, 1131177600, 1131181200, 1131184800, 
    1131188400, 1131192000, 1131195600, 1131199200, 1131202800, 1131206400, 
    1131210000, 1131213600, 1131217200, 1131220800, 1131224400, 1131228000, 
    1131231600, 1131235200, 1131238800, 1131242400, 1131246000, 1131249600, 
    1131253200, 1131256800, 1131260400, 1131264000, 1131267600, 1131271200, 
    1131274800, 1131278400, 1131282000, 1131285600, 1131289200, 1131292800, 
    1131296400, 1131300000, 1131303600, 1131307200, 1131310800, 1131314400, 
    1131318000, 1131321600, 1131325200, 1131328800, 1131332400, 1131336000, 
    1131339600, 1131343200, 1131346800, 1131350400, 1131354000, 1131357600, 
    1131361200, 1131364800, 1131368400, 1131372000, 1131375600, 1131379200, 
    1131382800, 1131386400, 1131390000, 1131393600, 1131397200, 1131400800, 
    1131404400, 1131408000, 1131411600, 1131415200, 1131418800, 1131422400, 
    1131426000, 1131429600, 1131433200, 1131436800, 1131440400, 1131444000, 
    1131447600, 1131451200, 1131454800, 1131458400, 1131462000, 1131465600, 
    1131469200, 1131472800, 1131476400, 1131480000, 1131483600, 1131487200, 
    1131490800, 1131494400, 1131498000, 1131501600, 1131505200, 1131508800, 
    1131512400, 1131516000, 1131519600, 1131523200, 1131526800, 1131530400, 
    1131534000, 1131537600, 1131541200, 1131544800, 1131548400, 1131552000, 
    1131555600, 1131559200, 1131562800, 1131566400, 1131570000, 1131573600, 
    1131577200, 1131580800, 1131584400, 1131588000, 1131591600, 1131595200, 
    1131598800, 1131602400, 1131606000, 1131609600, 1131613200, 1131616800, 
    1131620400, 1131624000, 1131627600, 1131631200, 1131634800, 1131638400, 
    1131642000, 1131645600, 1131649200, 1131652800, 1131656400, 1131660000, 
    1131663600, 1131667200, 1131670800, 1131674400, 1131678000, 1131681600, 
    1131685200, 1131688800, 1131692400, 1131696000, 1131699600, 1131703200, 
    1131706800, 1131710400, 1131714000, 1131717600, 1131721200, 1131724800, 
    1131728400, 1131732000, 1131735600, 1131739200, 1131742800, 1131746400, 
    1131750000, 1131753600, 1131757200, 1131760800, 1131764400, 1131768000, 
    1131771600, 1131775200, 1131778800, 1131782400, 1131786000, 1131789600, 
    1131793200, 1131796800, 1131800400, 1131804000, 1131807600, 1131811200, 
    1131814800, 1131818400, 1131822000, 1131825600, 1131829200, 1131832800, 
    1131836400, 1131840000, 1131843600, 1131847200, 1131850800, 1131854400, 
    1131858000, 1131861600, 1131865200, 1131868800, 1131872400, 1131876000, 
    1131879600, 1131883200, 1131886800, 1131890400, 1131894000, 1131897600, 
    1131901200, 1131904800, 1131908400, 1131912000, 1131915600, 1131919200, 
    1131922800, 1131926400, 1131930000, 1131933600, 1131937200, 1131940800, 
    1131944400, 1131948000, 1131951600, 1131955200, 1131958800, 1131962400, 
    1131966000, 1131969600, 1131973200, 1131976800, 1131980400, 1131984000, 
    1131987600, 1131991200, 1131994800, 1131998400, 1132002000, 1132005600, 
    1132009200, 1132012800, 1132016400, 1132020000, 1132023600, 1132027200, 
    1132030800, 1132034400, 1132038000, 1132041600, 1132045200, 1132048800, 
    1132052400, 1132056000, 1132059600, 1132063200, 1132066800, 1132070400, 
    1132074000, 1132077600, 1132081200, 1132084800, 1132088400, 1132092000, 
    1132095600, 1132099200, 1132102800, 1132106400, 1132110000, 1132113600, 
    1132117200, 1132120800, 1132124400, 1132128000, 1132131600, 1132135200, 
    1132138800, 1132142400, 1132146000, 1132149600, 1132153200, 1132156800, 
    1132160400, 1132164000, 1132167600, 1132171200, 1132174800, 1132178400, 
    1132182000, 1132185600, 1132189200, 1132192800, 1132196400, 1132200000, 
    1132203600, 1132207200, 1132210800, 1132214400, 1132218000, 1132221600, 
    1132225200, 1132228800, 1132232400, 1132236000, 1132239600, 1132243200, 
    1132246800, 1132250400, 1132254000, 1132257600, 1132261200, 1132264800, 
    1132268400, 1132272000, 1132275600, 1132279200, 1132282800, 1132286400, 
    1132290000, 1132293600, 1132297200, 1132300800, 1132304400, 1132308000, 
    1132311600, 1132315200, 1132318800, 1132322400, 1132326000, 1132329600, 
    1132333200, 1132336800, 1132340400, 1132344000, 1132347600, 1132351200, 
    1132354800, 1132358400, 1132362000, 1132365600, 1132369200, 1132372800, 
    1132376400, 1132380000, 1132383600, 1132387200, 1132390800, 1132394400, 
    1132398000, 1132401600, 1132405200, 1132408800, 1132412400, 1132416000, 
    1132419600, 1132423200, 1132426800, 1132430400, 1132434000, 1132437600, 
    1132441200, 1132444800, 1132448400, 1132452000, 1132455600, 1132459200, 
    1132462800, 1132466400, 1132470000, 1132473600, 1132477200, 1132480800, 
    1132484400, 1132488000, 1132491600, 1132495200, 1132498800, 1132502400, 
    1132506000, 1132509600, 1132513200, 1132516800, 1132520400, 1132524000, 
    1132527600, 1132531200, 1132534800, 1132538400, 1132542000, 1132545600, 
    1132549200, 1132552800, 1132556400, 1132560000, 1132563600, 1132567200, 
    1132570800, 1132574400, 1132578000, 1132581600, 1132585200, 1132588800, 
    1132592400, 1132596000, 1132599600, 1132603200, 1132606800, 1132610400, 
    1132614000, 1132617600, 1132621200, 1132624800, 1132628400, 1132632000, 
    1132635600, 1132639200, 1132642800, 1132646400, 1132650000, 1132653600, 
    1132657200, 1132660800, 1132664400, 1132668000, 1132671600, 1132675200, 
    1132678800, 1132682400, 1132686000, 1132689600, 1132693200, 1132696800, 
    1132700400, 1132704000, 1132707600, 1132711200, 1132714800, 1132718400, 
    1132722000, 1132725600, 1132729200, 1132732800, 1132736400, 1132740000, 
    1132743600, 1132747200, 1132750800, 1132754400, 1132758000, 1132761600, 
    1132765200, 1132768800, 1132772400, 1132776000, 1132779600, 1132783200, 
    1132786800, 1132790400, 1132794000, 1132797600, 1132801200, 1132804800, 
    1132808400, 1132812000, 1132815600, 1132819200, 1132822800, 1132826400, 
    1132830000, 1132833600, 1132837200, 1132840800, 1132844400, 1132848000, 
    1132851600, 1132855200, 1132858800, 1132862400, 1132866000, 1132869600, 
    1132873200, 1132876800, 1132880400, 1132884000, 1132887600, 1132891200, 
    1132894800, 1132898400, 1132902000, 1132905600, 1132909200, 1132912800, 
    1132916400, 1132920000, 1132923600, 1132927200, 1132930800, 1132934400, 
    1132938000, 1132941600, 1132945200, 1132948800, 1132952400, 1132956000, 
    1132959600, 1132963200, 1132966800, 1132970400, 1132974000, 1132977600, 
    1132981200, 1132984800, 1132988400, 1132992000, 1132995600, 1132999200, 
    1133002800, 1133006400, 1133010000, 1133013600, 1133017200, 1133020800, 
    1133024400, 1133028000, 1133031600, 1133035200, 1133038800, 1133042400, 
    1133046000, 1133049600, 1133053200, 1133056800, 1133060400, 1133064000, 
    1133067600, 1133071200, 1133074800, 1133078400, 1133082000, 1133085600, 
    1133089200, 1133092800, 1133096400, 1133100000, 1133103600, 1133107200, 
    1133110800, 1133114400, 1133118000, 1133121600, 1133125200, 1133128800, 
    1133132400, 1133136000, 1133139600, 1133143200, 1133146800, 1133150400, 
    1133154000, 1133157600, 1133161200, 1133164800, 1133168400, 1133172000, 
    1133175600, 1133179200, 1133182800, 1133186400, 1133190000, 1133193600, 
    1133197200, 1133200800, 1133204400, 1133208000, 1133211600, 1133215200, 
    1133218800, 1133222400, 1133226000, 1133229600, 1133233200, 1133236800, 
    1133240400, 1133244000, 1133247600, 1133251200, 1133254800, 1133258400, 
    1133262000, 1133265600, 1133269200, 1133272800, 1133276400, 1133280000, 
    1133283600, 1133287200, 1133290800, 1133294400, 1133298000, 1133301600, 
    1133305200, 1133308800, 1133312400, 1133316000, 1133319600, 1133323200, 
    1133326800, 1133330400, 1133334000, 1133337600, 1133341200, 1133344800, 
    1133348400, 1133352000, 1133355600, 1133359200, 1133362800, 1133366400, 
    1133370000, 1133373600, 1133377200, 1133380800, 1133384400, 1133388000, 
    1133391600, 1133395200, 1133398800, 1133402400, 1133406000, 1133409600, 
    1133413200, 1133416800, 1133420400, 1133424000, 1133427600, 1133431200, 
    1133434800, 1133438400, 1133442000, 1133445600, 1133449200, 1133452800, 
    1133456400, 1133460000, 1133463600, 1133467200, 1133470800, 1133474400, 
    1133478000, 1133481600, 1133485200, 1133488800, 1133492400, 1133496000, 
    1133499600, 1133503200, 1133506800, 1133510400, 1133514000, 1133517600, 
    1133521200, 1133524800, 1133528400, 1133532000, 1133535600, 1133539200, 
    1133542800, 1133546400, 1133550000, 1133553600, 1133557200, 1133560800, 
    1133564400, 1133568000, 1133571600, 1133575200, 1133578800, 1133582400, 
    1133586000, 1133589600, 1133593200, 1133596800, 1133600400, 1133604000, 
    1133607600, 1133611200, 1133614800, 1133618400, 1133622000, 1133625600, 
    1133629200, 1133632800, 1133636400, 1133640000, 1133643600, 1133647200, 
    1133650800, 1133654400, 1133658000, 1133661600, 1133665200, 1133668800, 
    1133672400, 1133676000, 1133679600, 1133683200, 1133686800, 1133690400, 
    1133694000, 1133697600, 1133701200, 1133704800, 1133708400, 1133712000, 
    1133715600, 1133719200, 1133722800, 1133726400, 1133730000, 1133733600, 
    1133737200, 1133740800, 1133744400, 1133748000, 1133751600, 1133755200, 
    1133758800, 1133762400, 1133766000, 1133769600, 1133773200, 1133776800, 
    1133780400, 1133784000, 1133787600, 1133791200, 1133794800, 1133798400, 
    1133802000, 1133805600, 1133809200, 1133812800, 1133816400, 1133820000, 
    1133823600, 1133827200, 1133830800, 1133834400, 1133838000, 1133841600, 
    1133845200, 1133848800, 1133852400, 1133856000, 1133859600, 1133863200, 
    1133866800, 1133870400, 1133874000, 1133877600, 1133881200, 1133884800, 
    1133888400, 1133892000, 1133895600, 1133899200, 1133902800, 1133906400, 
    1133910000, 1133913600, 1133917200, 1133920800, 1133924400, 1133928000, 
    1133931600, 1133935200, 1133938800, 1133942400, 1133946000, 1133949600, 
    1133953200, 1133956800, 1133960400, 1133964000, 1133967600, 1133971200, 
    1133974800, 1133978400, 1133982000, 1133985600, 1133989200, 1133992800, 
    1133996400, 1134000000, 1134003600, 1134007200, 1134010800, 1134014400, 
    1134018000, 1134021600, 1134025200, 1134028800, 1134032400, 1134036000, 
    1134039600, 1134043200, 1134046800, 1134050400, 1134054000, 1134057600, 
    1134061200, 1134064800, 1134068400, 1134072000, 1134075600, 1134079200, 
    1134082800, 1134086400, 1134090000, 1134093600, 1134097200, 1134100800, 
    1134104400, 1134108000, 1134111600, 1134115200, 1134118800, 1134122400, 
    1134126000, 1134129600, 1134133200, 1134136800, 1134140400, 1134144000, 
    1134147600, 1134151200, 1134154800, 1134158400, 1134162000, 1134165600, 
    1134169200, 1134172800, 1134176400, 1134180000, 1134183600, 1134187200, 
    1134190800, 1134194400, 1134198000, 1134201600, 1134205200, 1134208800, 
    1134212400, 1134216000, 1134219600, 1134223200, 1134226800, 1134230400, 
    1134234000, 1134237600, 1134241200, 1134244800, 1134248400, 1134252000, 
    1134255600, 1134259200, 1134262800, 1134266400, 1134270000, 1134273600, 
    1134277200, 1134280800, 1134284400, 1134288000, 1134291600, 1134295200, 
    1134298800, 1134302400, 1134306000, 1134309600, 1134313200, 1134316800, 
    1134320400, 1134324000, 1134327600, 1134331200, 1134334800, 1134338400, 
    1134342000, 1134345600, 1134349200, 1134352800, 1134356400, 1134360000, 
    1134363600, 1134367200, 1134370800, 1134374400, 1134378000, 1134381600, 
    1134385200, 1134388800, 1134392400, 1134396000, 1134399600, 1134403200, 
    1134406800, 1134410400, 1134414000, 1134417600, 1134421200, 1134424800, 
    1134428400, 1134432000, 1134435600, 1134439200, 1134442800, 1134446400, 
    1134450000, 1134453600, 1134457200, 1134460800, 1134464400, 1134468000, 
    1134471600, 1134475200, 1134478800, 1134482400, 1134486000, 1134489600, 
    1134493200, 1134496800, 1134500400, 1134504000, 1134507600, 1134511200, 
    1134514800, 1134518400, 1134522000, 1134525600, 1134529200, 1134532800, 
    1134536400, 1134540000, 1134543600, 1134547200, 1134550800, 1134554400, 
    1134558000, 1134561600, 1134565200, 1134568800, 1134572400, 1134576000, 
    1134579600, 1134583200, 1134586800, 1134590400, 1134594000, 1134597600, 
    1134601200, 1134604800, 1134608400, 1134612000, 1134615600, 1134619200, 
    1134622800, 1134626400, 1134630000, 1134633600, 1134637200, 1134640800, 
    1134644400, 1134648000, 1134651600, 1134655200, 1134658800, 1134662400, 
    1134666000, 1134669600, 1134673200, 1134676800, 1134680400, 1134684000, 
    1134687600, 1134691200, 1134694800, 1134698400, 1134702000, 1134705600, 
    1134709200, 1134712800, 1134716400, 1134720000, 1134723600, 1134727200, 
    1134730800, 1134734400, 1134738000, 1134741600, 1134745200, 1134748800, 
    1134752400, 1134756000, 1134759600, 1134763200, 1134766800, 1134770400, 
    1134774000, 1134777600, 1134781200, 1134784800, 1134788400, 1134792000, 
    1134795600, 1134799200, 1134802800, 1134806400, 1134810000, 1134813600, 
    1134817200, 1134820800, 1134824400, 1134828000, 1134831600, 1134835200, 
    1134838800, 1134842400, 1134846000, 1134849600, 1134853200, 1134856800, 
    1134860400, 1134864000, 1134867600, 1134871200, 1134874800, 1134878400, 
    1134882000, 1134885600, 1134889200, 1134892800, 1134896400, 1134900000, 
    1134903600, 1134907200, 1134910800, 1134914400, 1134918000, 1134921600, 
    1134925200, 1134928800, 1134932400, 1134936000, 1134939600, 1134943200, 
    1134946800, 1134950400, 1134954000, 1134957600, 1134961200, 1134964800, 
    1134968400, 1134972000, 1134975600, 1134979200, 1134982800, 1134986400, 
    1134990000, 1134993600, 1134997200, 1135000800, 1135004400, 1135008000, 
    1135011600, 1135015200, 1135018800, 1135022400, 1135026000, 1135029600, 
    1135033200, 1135036800, 1135040400, 1135044000, 1135047600, 1135051200, 
    1135054800, 1135058400, 1135062000, 1135065600, 1135069200, 1135072800, 
    1135076400, 1135080000, 1135083600, 1135087200, 1135090800, 1135094400, 
    1135098000, 1135101600, 1135105200, 1135108800, 1135112400, 1135116000, 
    1135119600, 1135123200, 1135126800, 1135130400, 1135134000, 1135137600, 
    1135141200, 1135144800, 1135148400, 1135152000, 1135155600, 1135159200, 
    1135162800, 1135166400, 1135170000, 1135173600, 1135177200, 1135180800, 
    1135184400, 1135188000, 1135191600, 1135195200, 1135198800, 1135202400, 
    1135206000, 1135209600, 1135213200, 1135216800, 1135220400, 1135224000, 
    1135227600, 1135231200, 1135234800, 1135238400, 1135242000, 1135245600, 
    1135249200, 1135252800, 1135256400, 1135260000, 1135263600, 1135267200, 
    1135270800, 1135274400, 1135278000, 1135281600, 1135285200, 1135288800, 
    1135292400, 1135296000, 1135299600, 1135303200, 1135306800, 1135310400, 
    1135314000, 1135317600, 1135321200, 1135324800, 1135328400, 1135332000, 
    1135335600, 1135339200, 1135342800, 1135346400, 1135350000, 1135353600, 
    1135357200, 1135360800, 1135364400, 1135368000, 1135371600, 1135375200, 
    1135378800, 1135382400, 1135386000, 1135389600, 1135393200, 1135396800, 
    1135400400, 1135404000, 1135407600, 1135411200, 1135414800, 1135418400, 
    1135422000, 1135425600, 1135429200, 1135432800, 1135436400, 1135440000, 
    1135443600, 1135447200, 1135450800, 1135454400, 1135458000, 1135461600, 
    1135465200, 1135468800, 1135472400, 1135476000, 1135479600, 1135483200, 
    1135486800, 1135490400, 1135494000, 1135497600, 1135501200, 1135504800, 
    1135508400, 1135512000, 1135515600, 1135519200, 1135522800, 1135526400, 
    1135530000, 1135533600, 1135537200, 1135540800, 1135544400, 1135548000, 
    1135551600, 1135555200, 1135558800, 1135562400, 1135566000, 1135569600, 
    1135573200, 1135576800, 1135580400, 1135584000, 1135587600, 1135591200, 
    1135594800, 1135598400, 1135602000, 1135605600, 1135609200, 1135612800, 
    1135616400, 1135620000, 1135623600, 1135627200, 1135630800, 1135634400, 
    1135638000, 1135641600, 1135645200, 1135648800, 1135652400, 1135656000, 
    1135659600, 1135663200, 1135666800, 1135670400, 1135674000, 1135677600, 
    1135681200, 1135684800, 1135688400, 1135692000, 1135695600, 1135699200, 
    1135702800, 1135706400, 1135710000, 1135713600, 1135717200, 1135720800, 
    1135724400, 1135728000, 1135731600, 1135735200, 1135738800, 1135742400, 
    1135746000, 1135749600, 1135753200, 1135756800, 1135760400, 1135764000, 
    1135767600, 1135771200, 1135774800, 1135778400, 1135782000, 1135785600, 
    1135789200, 1135792800, 1135796400, 1135800000, 1135803600, 1135807200, 
    1135810800, 1135814400, 1135818000, 1135821600, 1135825200, 1135828800, 
    1135832400, 1135836000, 1135839600, 1135843200, 1135846800, 1135850400, 
    1135854000, 1135857600, 1135861200, 1135864800, 1135868400, 1135872000, 
    1135875600, 1135879200, 1135882800, 1135886400, 1135890000, 1135893600, 
    1135897200, 1135900800, 1135904400, 1135908000, 1135911600, 1135915200, 
    1135918800, 1135922400, 1135926000, 1135929600, 1135933200, 1135936800, 
    1135940400, 1135944000, 1135947600, 1135951200, 1135954800, 1135958400, 
    1135962000, 1135965600, 1135969200, 1135972800, 1135976400, 1135980000, 
    1135983600, 1135987200, 1135990800, 1135994400, 1135998000, 1136001600, 
    1136005200, 1136008800, 1136012400, 1136016000, 1136019600, 1136023200, 
    1136026800, 1136030400, 1136034000, 1136037600, 1136041200, 1136044800, 
    1136048400, 1136052000, 1136055600, 1136059200, 1136062800, 1136066400, 
    1136070000, 1136073600, 1136077200, 1136080800, 1136084400, 1136088000, 
    1136091600, 1136095200, 1136098800, 1136102400, 1136106000, 1136109600, 
    1136113200, 1136116800, 1136120400, 1136124000, 1136127600, 1136131200, 
    1136134800, 1136138400, 1136142000, 1136145600, 1136149200, 1136152800, 
    1136156400, 1136160000, 1136163600, 1136167200, 1136170800, 1136174400, 
    1136178000, 1136181600, 1136185200, 1136188800, 1136192400, 1136196000, 
    1136199600, 1136203200, 1136206800, 1136210400, 1136214000, 1136217600, 
    1136221200, 1136224800, 1136228400, 1136232000, 1136235600, 1136239200, 
    1136242800, 1136246400, 1136250000, 1136253600, 1136257200, 1136260800, 
    1136264400, 1136268000, 1136271600, 1136275200, 1136278800, 1136282400, 
    1136286000, 1136289600, 1136293200, 1136296800, 1136300400, 1136304000, 
    1136307600, 1136311200, 1136314800, 1136318400, 1136322000, 1136325600, 
    1136329200, 1136332800, 1136336400, 1136340000, 1136343600, 1136347200, 
    1136350800, 1136354400, 1136358000, 1136361600, 1136365200, 1136368800, 
    1136372400, 1136376000, 1136379600, 1136383200, 1136386800, 1136390400, 
    1136394000, 1136397600, 1136401200, 1136404800, 1136408400, 1136412000, 
    1136415600, 1136419200, 1136422800, 1136426400, 1136430000, 1136433600, 
    1136437200, 1136440800, 1136444400, 1136448000, 1136451600, 1136455200, 
    1136458800, 1136462400, 1136466000, 1136469600, 1136473200, 1136476800, 
    1136480400, 1136484000, 1136487600, 1136491200, 1136494800, 1136498400, 
    1136502000, 1136505600, 1136509200, 1136512800, 1136516400, 1136520000, 
    1136523600, 1136527200, 1136530800, 1136534400, 1136538000, 1136541600, 
    1136545200, 1136548800, 1136552400, 1136556000, 1136559600, 1136563200, 
    1136566800, 1136570400, 1136574000, 1136577600, 1136581200, 1136584800, 
    1136588400, 1136592000, 1136595600, 1136599200, 1136602800, 1136606400, 
    1136610000, 1136613600, 1136617200, 1136620800, 1136624400, 1136628000, 
    1136631600, 1136635200, 1136638800, 1136642400, 1136646000, 1136649600, 
    1136653200, 1136656800, 1136660400, 1136664000, 1136667600, 1136671200, 
    1136674800, 1136678400, 1136682000, 1136685600, 1136689200, 1136692800, 
    1136696400, 1136700000, 1136703600, 1136707200, 1136710800, 1136714400, 
    1136718000, 1136721600, 1136725200, 1136728800, 1136732400, 1136736000, 
    1136739600, 1136743200, 1136746800, 1136750400, 1136754000, 1136757600, 
    1136761200, 1136764800, 1136768400, 1136772000, 1136775600, 1136779200, 
    1136782800, 1136786400, 1136790000, 1136793600, 1136797200, 1136800800, 
    1136804400, 1136808000, 1136811600, 1136815200, 1136818800, 1136822400, 
    1136826000, 1136829600, 1136833200, 1136836800, 1136840400, 1136844000, 
    1136847600, 1136851200, 1136854800, 1136858400, 1136862000, 1136865600, 
    1136869200, 1136872800, 1136876400, 1136880000, 1136883600, 1136887200, 
    1136890800, 1136894400, 1136898000, 1136901600, 1136905200, 1136908800, 
    1136912400, 1136916000, 1136919600, 1136923200, 1136926800, 1136930400, 
    1136934000, 1136937600, 1136941200, 1136944800, 1136948400, 1136952000, 
    1136955600, 1136959200, 1136962800, 1136966400, 1136970000, 1136973600, 
    1136977200, 1136980800, 1136984400, 1136988000, 1136991600, 1136995200, 
    1136998800, 1137002400, 1137006000, 1137009600, 1137013200, 1137016800, 
    1137020400, 1137024000, 1137027600, 1137031200, 1137034800, 1137038400, 
    1137042000, 1137045600, 1137049200, 1137052800, 1137056400, 1137060000, 
    1137063600, 1137067200, 1137070800, 1137074400, 1137078000, 1137081600, 
    1137085200, 1137088800, 1137092400, 1137096000, 1137099600, 1137103200, 
    1137106800, 1137110400, 1137114000, 1137117600, 1137121200, 1137124800, 
    1137128400, 1137132000, 1137135600, 1137139200, 1137142800, 1137146400, 
    1137150000, 1137153600, 1137157200, 1137160800, 1137164400, 1137168000, 
    1137171600, 1137175200, 1137178800, 1137182400, 1137186000, 1137189600, 
    1137193200, 1137196800, 1137200400, 1137204000, 1137207600, 1137211200, 
    1137214800, 1137218400, 1137222000, 1137225600, 1137229200, 1137232800, 
    1137236400, 1137240000, 1137243600, 1137247200, 1137250800, 1137254400, 
    1137258000, 1137261600, 1137265200, 1137268800, 1137272400, 1137276000, 
    1137279600, 1137283200, 1137286800, 1137290400, 1137294000, 1137297600, 
    1137301200, 1137304800, 1137308400, 1137312000, 1137315600, 1137319200, 
    1137322800, 1137326400, 1137330000, 1137333600, 1137337200, 1137340800, 
    1137344400, 1137348000, 1137351600, 1137355200, 1137358800, 1137362400, 
    1137366000, 1137369600, 1137373200, 1137376800, 1137380400, 1137384000, 
    1137387600, 1137391200, 1137394800, 1137398400, 1137402000, 1137405600, 
    1137409200, 1137412800, 1137416400, 1137420000, 1137423600, 1137427200, 
    1137430800, 1137434400, 1137438000, 1137441600, 1137445200, 1137448800, 
    1137452400, 1137456000, 1137459600, 1137463200, 1137466800, 1137470400, 
    1137474000, 1137477600, 1137481200, 1137484800, 1137488400, 1137492000, 
    1137495600, 1137499200, 1137502800, 1137506400, 1137510000, 1137513600, 
    1137517200, 1137520800, 1137524400, 1137528000, 1137531600, 1137535200, 
    1137538800, 1137542400, 1137546000, 1137549600, 1137553200, 1137556800, 
    1137560400, 1137564000, 1137567600, 1137571200, 1137574800, 1137578400, 
    1137582000, 1137585600, 1137589200, 1137592800, 1137596400, 1137600000, 
    1137603600, 1137607200, 1137610800, 1137614400, 1137618000, 1137621600, 
    1137625200, 1137628800, 1137632400, 1137636000, 1137639600, 1137643200, 
    1137646800, 1137650400, 1137654000, 1137657600, 1137661200, 1137664800, 
    1137668400, 1137672000, 1137675600, 1137679200, 1137682800, 1137686400, 
    1137690000, 1137693600, 1137697200, 1137700800, 1137704400, 1137708000, 
    1137711600, 1137715200, 1137718800, 1137722400, 1137726000, 1137729600, 
    1137733200, 1137736800, 1137740400, 1137744000, 1137747600, 1137751200, 
    1137754800, 1137758400, 1137762000, 1137765600, 1137769200, 1137772800, 
    1137776400, 1137780000, 1137783600, 1137787200, 1137790800, 1137794400, 
    1137798000, 1137801600, 1137805200, 1137808800, 1137812400, 1137816000, 
    1137819600, 1137823200, 1137826800, 1137830400, 1137834000, 1137837600, 
    1137841200, 1137844800, 1137848400, 1137852000, 1137855600, 1137859200, 
    1137862800, 1137866400, 1137870000, 1137873600, 1137877200, 1137880800, 
    1137884400, 1137888000, 1137891600, 1137895200, 1137898800, 1137902400, 
    1137906000, 1137909600, 1137913200, 1137916800, 1137920400, 1137924000, 
    1137927600, 1137931200, 1137934800, 1137938400, 1137942000, 1137945600, 
    1137949200, 1137952800, 1137956400, 1137960000, 1137963600, 1137967200, 
    1137970800, 1137974400, 1137978000, 1137981600, 1137985200, 1137988800, 
    1137992400, 1137996000, 1137999600, 1138003200, 1138006800, 1138010400, 
    1138014000, 1138017600, 1138021200, 1138024800, 1138028400, 1138032000, 
    1138035600, 1138039200, 1138042800, 1138046400, 1138050000, 1138053600, 
    1138057200, 1138060800, 1138064400, 1138068000, 1138071600, 1138075200, 
    1138078800, 1138082400, 1138086000, 1138089600, 1138093200, 1138096800, 
    1138100400, 1138104000, 1138107600, 1138111200, 1138114800, 1138118400, 
    1138122000, 1138125600, 1138129200, 1138132800, 1138136400, 1138140000, 
    1138143600, 1138147200, 1138150800, 1138154400, 1138158000, 1138161600, 
    1138165200, 1138168800, 1138172400, 1138176000, 1138179600, 1138183200, 
    1138186800, 1138190400, 1138194000, 1138197600, 1138201200, 1138204800, 
    1138208400, 1138212000, 1138215600, 1138219200, 1138222800, 1138226400, 
    1138230000, 1138233600, 1138237200, 1138240800, 1138244400, 1138248000, 
    1138251600, 1138255200, 1138258800, 1138262400, 1138266000, 1138269600, 
    1138273200, 1138276800, 1138280400, 1138284000, 1138287600, 1138291200, 
    1138294800, 1138298400, 1138302000, 1138305600, 1138309200, 1138312800, 
    1138316400, 1138320000, 1138323600, 1138327200, 1138330800, 1138334400, 
    1138338000, 1138341600, 1138345200, 1138348800, 1138352400, 1138356000, 
    1138359600, 1138363200, 1138366800, 1138370400, 1138374000, 1138377600, 
    1138381200, 1138384800, 1138388400, 1138392000, 1138395600, 1138399200, 
    1138402800, 1138406400, 1138410000, 1138413600, 1138417200, 1138420800, 
    1138424400, 1138428000, 1138431600, 1138435200, 1138438800, 1138442400, 
    1138446000, 1138449600, 1138453200, 1138456800, 1138460400, 1138464000, 
    1138467600, 1138471200, 1138474800, 1138478400, 1138482000, 1138485600, 
    1138489200, 1138492800, 1138496400, 1138500000, 1138503600, 1138507200, 
    1138510800, 1138514400, 1138518000, 1138521600, 1138525200, 1138528800, 
    1138532400, 1138536000, 1138539600, 1138543200, 1138546800, 1138550400, 
    1138554000, 1138557600, 1138561200, 1138564800, 1138568400, 1138572000, 
    1138575600, 1138579200, 1138582800, 1138586400, 1138590000, 1138593600, 
    1138597200, 1138600800, 1138604400, 1138608000, 1138611600, 1138615200, 
    1138618800, 1138622400, 1138626000, 1138629600, 1138633200, 1138636800, 
    1138640400, 1138644000, 1138647600, 1138651200, 1138654800, 1138658400, 
    1138662000, 1138665600, 1138669200, 1138672800, 1138676400, 1138680000, 
    1138683600, 1138687200, 1138690800, 1138694400, 1138698000, 1138701600, 
    1138705200, 1138708800, 1138712400, 1138716000, 1138719600, 1138723200, 
    1138726800, 1138730400, 1138734000, 1138737600, 1138741200, 1138744800, 
    1138748400, 1138752000, 1138755600, 1138759200, 1138762800, 1138766400, 
    1138770000, 1138773600, 1138777200, 1138780800, 1138784400, 1138788000, 
    1138791600, 1138795200, 1138798800, 1138802400, 1138806000, 1138809600, 
    1138813200, 1138816800, 1138820400, 1138824000, 1138827600, 1138831200, 
    1138834800, 1138838400, 1138842000, 1138845600, 1138849200, 1138852800, 
    1138856400, 1138860000, 1138863600, 1138867200, 1138870800, 1138874400, 
    1138878000, 1138881600, 1138885200, 1138888800, 1138892400, 1138896000, 
    1138899600, 1138903200, 1138906800, 1138910400, 1138914000, 1138917600, 
    1138921200, 1138924800, 1138928400, 1138932000, 1138935600, 1138939200, 
    1138942800, 1138946400, 1138950000, 1138953600, 1138957200, 1138960800, 
    1138964400, 1138968000, 1138971600, 1138975200, 1138978800, 1138982400, 
    1138986000, 1138989600, 1138993200, 1138996800, 1139000400, 1139004000, 
    1139007600, 1139011200, 1139014800, 1139018400, 1139022000, 1139025600, 
    1139029200, 1139032800, 1139036400, 1139040000, 1139043600, 1139047200, 
    1139050800, 1139054400, 1139058000, 1139061600, 1139065200, 1139068800, 
    1139072400, 1139076000, 1139079600, 1139083200, 1139086800, 1139090400, 
    1139094000, 1139097600, 1139101200, 1139104800, 1139108400, 1139112000, 
    1139115600, 1139119200, 1139122800, 1139126400, 1139130000, 1139133600, 
    1139137200, 1139140800, 1139144400, 1139148000, 1139151600, 1139155200, 
    1139158800, 1139162400, 1139166000, 1139169600, 1139173200, 1139176800, 
    1139180400, 1139184000, 1139187600, 1139191200, 1139194800, 1139198400, 
    1139202000, 1139205600, 1139209200, 1139212800, 1139216400, 1139220000, 
    1139223600, 1139227200, 1139230800, 1139234400, 1139238000, 1139241600, 
    1139245200, 1139248800, 1139252400, 1139256000, 1139259600, 1139263200, 
    1139266800, 1139270400, 1139274000, 1139277600, 1139281200, 1139284800, 
    1139288400, 1139292000, 1139295600, 1139299200, 1139302800, 1139306400, 
    1139310000, 1139313600, 1139317200, 1139320800, 1139324400, 1139328000, 
    1139331600, 1139335200, 1139338800, 1139342400, 1139346000, 1139349600, 
    1139353200, 1139356800, 1139360400, 1139364000, 1139367600, 1139371200, 
    1139374800, 1139378400, 1139382000, 1139385600, 1139389200, 1139392800, 
    1139396400, 1139400000, 1139403600, 1139407200, 1139410800, 1139414400, 
    1139418000, 1139421600, 1139425200, 1139428800, 1139432400, 1139436000, 
    1139439600, 1139443200, 1139446800, 1139450400, 1139454000, 1139457600, 
    1139461200, 1139464800, 1139468400, 1139472000, 1139475600, 1139479200, 
    1139482800, 1139486400, 1139490000, 1139493600, 1139497200, 1139500800, 
    1139504400, 1139508000, 1139511600, 1139515200, 1139518800, 1139522400, 
    1139526000, 1139529600, 1139533200, 1139536800, 1139540400, 1139544000, 
    1139547600, 1139551200, 1139554800, 1139558400, 1139562000, 1139565600, 
    1139569200, 1139572800, 1139576400, 1139580000, 1139583600, 1139587200, 
    1139590800, 1139594400, 1139598000, 1139601600, 1139605200, 1139608800, 
    1139612400, 1139616000, 1139619600, 1139623200, 1139626800, 1139630400, 
    1139634000, 1139637600, 1139641200, 1139644800, 1139648400, 1139652000, 
    1139655600, 1139659200, 1139662800, 1139666400, 1139670000, 1139673600, 
    1139677200, 1139680800, 1139684400, 1139688000, 1139691600, 1139695200, 
    1139698800, 1139702400, 1139706000, 1139709600, 1139713200, 1139716800, 
    1139720400, 1139724000, 1139727600, 1139731200, 1139734800, 1139738400, 
    1139742000, 1139745600, 1139749200, 1139752800, 1139756400, 1139760000, 
    1139763600, 1139767200, 1139770800, 1139774400, 1139778000, 1139781600, 
    1139785200, 1139788800, 1139792400, 1139796000, 1139799600, 1139803200, 
    1139806800, 1139810400, 1139814000, 1139817600, 1139821200, 1139824800, 
    1139828400, 1139832000, 1139835600, 1139839200, 1139842800, 1139846400, 
    1139850000, 1139853600, 1139857200, 1139860800, 1139864400, 1139868000, 
    1139871600, 1139875200, 1139878800, 1139882400, 1139886000, 1139889600, 
    1139893200, 1139896800, 1139900400, 1139904000, 1139907600, 1139911200, 
    1139914800, 1139918400, 1139922000, 1139925600, 1139929200, 1139932800, 
    1139936400, 1139940000, 1139943600, 1139947200, 1139950800, 1139954400, 
    1139958000, 1139961600, 1139965200, 1139968800, 1139972400, 1139976000, 
    1139979600, 1139983200, 1139986800, 1139990400, 1139994000, 1139997600, 
    1140001200, 1140004800, 1140008400, 1140012000, 1140015600, 1140019200, 
    1140022800, 1140026400, 1140030000, 1140033600, 1140037200, 1140040800, 
    1140044400, 1140048000, 1140051600, 1140055200, 1140058800, 1140062400, 
    1140066000, 1140069600, 1140073200, 1140076800, 1140080400, 1140084000, 
    1140087600, 1140091200, 1140094800, 1140098400, 1140102000, 1140105600, 
    1140109200, 1140112800, 1140116400, 1140120000, 1140123600, 1140127200, 
    1140130800, 1140134400, 1140138000, 1140141600, 1140145200, 1140148800, 
    1140152400, 1140156000, 1140159600, 1140163200, 1140166800, 1140170400, 
    1140174000, 1140177600, 1140181200, 1140184800, 1140188400, 1140192000, 
    1140195600, 1140199200, 1140202800, 1140206400, 1140210000, 1140213600, 
    1140217200, 1140220800, 1140224400, 1140228000, 1140231600, 1140235200, 
    1140238800, 1140242400, 1140246000, 1140249600, 1140253200, 1140256800, 
    1140260400, 1140264000, 1140267600, 1140271200, 1140274800, 1140278400, 
    1140282000, 1140285600, 1140289200, 1140292800, 1140296400, 1140300000, 
    1140303600, 1140307200, 1140310800, 1140314400, 1140318000, 1140321600, 
    1140325200, 1140328800, 1140332400, 1140336000, 1140339600, 1140343200, 
    1140346800, 1140350400, 1140354000, 1140357600, 1140361200, 1140364800, 
    1140368400, 1140372000, 1140375600, 1140379200, 1140382800, 1140386400, 
    1140390000, 1140393600, 1140397200, 1140400800, 1140404400, 1140408000, 
    1140411600, 1140415200, 1140418800, 1140422400, 1140426000, 1140429600, 
    1140433200, 1140436800, 1140440400, 1140444000, 1140447600, 1140451200, 
    1140454800, 1140458400, 1140462000, 1140465600, 1140469200, 1140472800, 
    1140476400, 1140480000, 1140483600, 1140487200, 1140490800, 1140494400, 
    1140498000, 1140501600, 1140505200, 1140508800, 1140512400, 1140516000, 
    1140519600, 1140523200, 1140526800, 1140530400, 1140534000, 1140537600, 
    1140541200, 1140544800, 1140548400, 1140552000, 1140555600, 1140559200, 
    1140562800, 1140566400, 1140570000, 1140573600, 1140577200, 1140580800, 
    1140584400, 1140588000, 1140591600, 1140595200, 1140598800, 1140602400, 
    1140606000, 1140609600, 1140613200, 1140616800, 1140620400, 1140624000, 
    1140627600, 1140631200, 1140634800, 1140638400, 1140642000, 1140645600, 
    1140649200, 1140652800, 1140656400, 1140660000, 1140663600, 1140667200, 
    1140670800, 1140674400, 1140678000, 1140681600, 1140685200, 1140688800, 
    1140692400, 1140696000, 1140699600, 1140703200, 1140706800, 1140710400, 
    1140714000, 1140717600, 1140721200, 1140724800, 1140728400, 1140732000, 
    1140735600, 1140739200, 1140742800, 1140746400, 1140750000, 1140753600, 
    1140757200, 1140760800, 1140764400, 1140768000, 1140771600, 1140775200, 
    1140778800, 1140782400, 1140786000, 1140789600, 1140793200, 1140796800, 
    1140800400, 1140804000, 1140807600, 1140811200, 1140814800, 1140818400, 
    1140822000, 1140825600, 1140829200, 1140832800, 1140836400, 1140840000, 
    1140843600, 1140847200, 1140850800, 1140854400, 1140858000, 1140861600, 
    1140865200, 1140868800, 1140872400, 1140876000, 1140879600, 1140883200, 
    1140886800, 1140890400, 1140894000, 1140897600, 1140901200, 1140904800, 
    1140908400, 1140912000, 1140915600, 1140919200, 1140922800, 1140926400, 
    1140930000, 1140933600, 1140937200, 1140940800, 1140944400, 1140948000, 
    1140951600, 1140955200, 1140958800, 1140962400, 1140966000, 1140969600, 
    1140973200, 1140976800, 1140980400, 1140984000, 1140987600, 1140991200, 
    1140994800, 1140998400, 1141002000, 1141005600, 1141009200, 1141012800, 
    1141016400, 1141020000, 1141023600, 1141027200, 1141030800, 1141034400, 
    1141038000, 1141041600, 1141045200, 1141048800, 1141052400, 1141056000, 
    1141059600, 1141063200, 1141066800, 1141070400, 1141074000, 1141077600, 
    1141081200, 1141084800, 1141088400, 1141092000, 1141095600, 1141099200, 
    1141102800, 1141106400, 1141110000, 1141113600, 1141117200, 1141120800, 
    1141124400, 1141128000, 1141131600, 1141135200, 1141138800, 1141142400, 
    1141146000, 1141149600, 1141153200, 1141156800, 1141160400, 1141164000, 
    1141167600, 1141171200, 1141174800, 1141178400, 1141182000, 1141185600, 
    1141189200, 1141192800, 1141196400, 1141200000, 1141203600, 1141207200, 
    1141210800, 1141214400, 1141218000, 1141221600, 1141225200, 1141228800, 
    1141232400, 1141236000, 1141239600, 1141243200, 1141246800, 1141250400, 
    1141254000, 1141257600, 1141261200, 1141264800, 1141268400, 1141272000, 
    1141275600, 1141279200, 1141282800, 1141286400, 1141290000, 1141293600, 
    1141297200, 1141300800, 1141304400, 1141308000, 1141311600, 1141315200, 
    1141318800, 1141322400, 1141326000, 1141329600, 1141333200, 1141336800, 
    1141340400, 1141344000, 1141347600, 1141351200, 1141354800, 1141358400, 
    1141362000, 1141365600, 1141369200, 1141372800, 1141376400, 1141380000, 
    1141383600, 1141387200, 1141390800, 1141394400, 1141398000, 1141401600, 
    1141405200, 1141408800, 1141412400, 1141416000, 1141419600, 1141423200, 
    1141426800, 1141430400, 1141434000, 1141437600, 1141441200, 1141444800, 
    1141448400, 1141452000, 1141455600, 1141459200, 1141462800, 1141466400, 
    1141470000, 1141473600, 1141477200, 1141480800, 1141484400, 1141488000, 
    1141491600, 1141495200, 1141498800, 1141502400, 1141506000, 1141509600, 
    1141513200, 1141516800, 1141520400, 1141524000, 1141527600, 1141531200, 
    1141534800, 1141538400, 1141542000, 1141545600, 1141549200, 1141552800, 
    1141556400, 1141560000, 1141563600, 1141567200, 1141570800, 1141574400, 
    1141578000, 1141581600, 1141585200, 1141588800, 1141592400, 1141596000, 
    1141599600, 1141603200, 1141606800, 1141610400, 1141614000, 1141617600, 
    1141621200, 1141624800, 1141628400, 1141632000, 1141635600, 1141639200, 
    1141642800, 1141646400, 1141650000, 1141653600, 1141657200, 1141660800, 
    1141664400, 1141668000, 1141671600, 1141675200, 1141678800, 1141682400, 
    1141686000, 1141689600, 1141693200, 1141696800, 1141700400, 1141704000, 
    1141707600, 1141711200, 1141714800, 1141718400, 1141722000, 1141725600, 
    1141729200, 1141732800, 1141736400, 1141740000, 1141743600, 1141747200, 
    1141750800, 1141754400, 1141758000, 1141761600, 1141765200, 1141768800, 
    1141772400, 1141776000, 1141779600, 1141783200, 1141786800, 1141790400, 
    1141794000, 1141797600, 1141801200, 1141804800, 1141808400, 1141812000, 
    1141815600, 1141819200, 1141822800, 1141826400, 1141830000, 1141833600, 
    1141837200, 1141840800, 1141844400, 1141848000, 1141851600, 1141855200, 
    1141858800, 1141862400, 1141866000, 1141869600, 1141873200, 1141876800, 
    1141880400, 1141884000, 1141887600, 1141891200, 1141894800, 1141898400, 
    1141902000, 1141905600, 1141909200, 1141912800, 1141916400, 1141920000, 
    1141923600, 1141927200, 1141930800, 1141934400, 1141938000, 1141941600, 
    1141945200, 1141948800, 1141952400, 1141956000, 1141959600, 1141963200, 
    1141966800, 1141970400, 1141974000, 1141977600, 1141981200, 1141984800, 
    1141988400, 1141992000, 1141995600, 1141999200, 1142002800, 1142006400, 
    1142010000, 1142013600, 1142017200, 1142020800, 1142024400, 1142028000, 
    1142031600, 1142035200, 1142038800, 1142042400, 1142046000, 1142049600, 
    1142053200, 1142056800, 1142060400, 1142064000, 1142067600, 1142071200, 
    1142074800, 1142078400, 1142082000, 1142085600, 1142089200, 1142092800, 
    1142096400, 1142100000, 1142103600, 1142107200, 1142110800, 1142114400, 
    1142118000, 1142121600, 1142125200, 1142128800, 1142132400, 1142136000, 
    1142139600, 1142143200, 1142146800, 1142150400, 1142154000, 1142157600, 
    1142161200, 1142164800, 1142168400, 1142172000, 1142175600, 1142179200, 
    1142182800, 1142186400, 1142190000, 1142193600, 1142197200, 1142200800, 
    1142204400, 1142208000, 1142211600, 1142215200, 1142218800, 1142222400, 
    1142226000, 1142229600, 1142233200, 1142236800, 1142240400, 1142244000, 
    1142247600, 1142251200, 1142254800, 1142258400, 1142262000, 1142265600, 
    1142269200, 1142272800, 1142276400, 1142280000, 1142283600, 1142287200, 
    1142290800, 1142294400, 1142298000, 1142301600, 1142305200, 1142308800, 
    1142312400, 1142316000, 1142319600, 1142323200, 1142326800, 1142330400, 
    1142334000, 1142337600, 1142341200, 1142344800, 1142348400, 1142352000, 
    1142355600, 1142359200, 1142362800, 1142366400, 1142370000, 1142373600, 
    1142377200, 1142380800, 1142384400, 1142388000, 1142391600, 1142395200, 
    1142398800, 1142402400, 1142406000, 1142409600, 1142413200, 1142416800, 
    1142420400, 1142424000, 1142427600, 1142431200, 1142434800, 1142438400, 
    1142442000, 1142445600, 1142449200, 1142452800, 1142456400, 1142460000, 
    1142463600, 1142467200, 1142470800, 1142474400, 1142478000, 1142481600, 
    1142485200, 1142488800, 1142492400, 1142496000, 1142499600, 1142503200, 
    1142506800, 1142510400, 1142514000, 1142517600, 1142521200, 1142524800, 
    1142528400, 1142532000, 1142535600, 1142539200, 1142542800, 1142546400, 
    1142550000, 1142553600, 1142557200, 1142560800, 1142564400, 1142568000, 
    1142571600, 1142575200, 1142578800, 1142582400, 1142586000, 1142589600, 
    1142593200, 1142596800, 1142600400, 1142604000, 1142607600, 1142611200, 
    1142614800, 1142618400, 1142622000, 1142625600, 1142629200, 1142632800, 
    1142636400, 1142640000, 1142643600, 1142647200, 1142650800, 1142654400, 
    1142658000, 1142661600, 1142665200, 1142668800, 1142672400, 1142676000, 
    1142679600, 1142683200, 1142686800, 1142690400, 1142694000, 1142697600, 
    1142701200, 1142704800, 1142708400, 1142712000, 1142715600, 1142719200, 
    1142722800, 1142726400, 1142730000, 1142733600, 1142737200, 1142740800, 
    1142744400, 1142748000, 1142751600, 1142755200, 1142758800, 1142762400, 
    1142766000, 1142769600, 1142773200, 1142776800, 1142780400, 1142784000, 
    1142787600, 1142791200, 1142794800, 1142798400, 1142802000, 1142805600, 
    1142809200, 1142812800, 1142816400, 1142820000, 1142823600, 1142827200, 
    1142830800, 1142834400, 1142838000, 1142841600, 1142845200, 1142848800, 
    1142852400, 1142856000, 1142859600, 1142863200, 1142866800, 1142870400, 
    1142874000, 1142877600, 1142881200, 1142884800, 1142888400, 1142892000, 
    1142895600, 1142899200, 1142902800, 1142906400, 1142910000, 1142913600, 
    1142917200, 1142920800, 1142924400, 1142928000, 1142931600, 1142935200, 
    1142938800, 1142942400, 1142946000, 1142949600, 1142953200, 1142956800, 
    1142960400, 1142964000, 1142967600, 1142971200, 1142974800, 1142978400, 
    1142982000, 1142985600, 1142989200, 1142992800, 1142996400, 1143000000, 
    1143003600, 1143007200, 1143010800, 1143014400, 1143018000, 1143021600, 
    1143025200, 1143028800, 1143032400, 1143036000, 1143039600, 1143043200, 
    1143046800, 1143050400, 1143054000, 1143057600, 1143061200, 1143064800, 
    1143068400, 1143072000, 1143075600, 1143079200, 1143082800, 1143086400, 
    1143090000, 1143093600, 1143097200, 1143100800, 1143104400, 1143108000, 
    1143111600, 1143115200, 1143118800, 1143122400, 1143126000, 1143129600, 
    1143133200, 1143136800, 1143140400, 1143144000, 1143147600, 1143151200, 
    1143154800, 1143158400, 1143162000, 1143165600, 1143169200, 1143172800, 
    1143176400, 1143180000, 1143183600, 1143187200, 1143190800, 1143194400, 
    1143198000, 1143201600, 1143205200, 1143208800, 1143212400, 1143216000, 
    1143219600, 1143223200, 1143226800, 1143230400, 1143234000, 1143237600, 
    1143241200, 1143244800, 1143248400, 1143252000, 1143255600, 1143259200, 
    1143262800, 1143266400, 1143270000, 1143273600, 1143277200, 1143280800, 
    1143284400, 1143288000, 1143291600, 1143295200, 1143298800, 1143302400, 
    1143306000, 1143309600, 1143313200, 1143316800, 1143320400, 1143324000, 
    1143327600, 1143331200, 1143334800, 1143338400, 1143342000, 1143345600, 
    1143349200, 1143352800, 1143356400, 1143360000, 1143363600, 1143367200, 
    1143370800, 1143374400, 1143378000, 1143381600, 1143385200, 1143388800, 
    1143392400, 1143396000, 1143399600, 1143403200, 1143406800, 1143410400, 
    1143414000, 1143417600, 1143421200, 1143424800, 1143428400, 1143432000, 
    1143435600, 1143439200, 1143442800, 1143446400, 1143450000, 1143453600, 
    1143457200, 1143460800, 1143464400, 1143468000, 1143471600, 1143475200, 
    1143478800, 1143482400, 1143486000, 1143489600, 1143493200, 1143496800, 
    1143500400, 1143504000, 1143507600, 1143511200, 1143514800, 1143518400, 
    1143522000, 1143525600, 1143529200, 1143532800, 1143536400, 1143540000, 
    1143543600, 1143547200, 1143550800, 1143554400, 1143558000, 1143561600, 
    1143565200, 1143568800, 1143572400, 1143576000, 1143579600, 1143583200, 
    1143586800, 1143590400, 1143594000, 1143597600, 1143601200, 1143604800, 
    1143608400, 1143612000, 1143615600, 1143619200, 1143622800, 1143626400, 
    1143630000, 1143633600, 1143637200, 1143640800, 1143644400, 1143648000, 
    1143651600, 1143655200, 1143658800, 1143662400, 1143666000, 1143669600, 
    1143673200, 1143676800, 1143680400, 1143684000, 1143687600, 1143691200, 
    1143694800, 1143698400, 1143702000, 1143705600, 1143709200, 1143712800, 
    1143716400, 1143720000, 1143723600, 1143727200, 1143730800, 1143734400, 
    1143738000, 1143741600, 1143745200, 1143748800, 1143752400, 1143756000, 
    1143759600, 1143763200, 1143766800, 1143770400, 1143774000, 1143777600, 
    1143781200, 1143784800, 1143788400, 1143792000, 1143795600, 1143799200, 
    1143802800, 1143806400, 1143810000, 1143813600, 1143817200, 1143820800, 
    1143824400, 1143828000, 1143831600, 1143835200, 1143838800, 1143842400, 
    1143846000, 1143849600, 1143853200, 1143856800, 1143860400, 1143864000, 
    1143867600, 1143871200, 1143874800, 1143878400, 1143882000, 1143885600, 
    1143889200, 1143892800, 1143896400, 1143900000, 1143903600, 1143907200, 
    1143910800, 1143914400, 1143918000, 1143921600, 1143925200, 1143928800, 
    1143932400, 1143936000, 1143939600, 1143943200, 1143946800, 1143950400, 
    1143954000, 1143957600, 1143961200, 1143964800, 1143968400, 1143972000, 
    1143975600, 1143979200, 1143982800, 1143986400, 1143990000, 1143993600, 
    1143997200, 1144000800, 1144004400, 1144008000, 1144011600, 1144015200, 
    1144018800, 1144022400, 1144026000, 1144029600, 1144033200, 1144036800, 
    1144040400, 1144044000, 1144047600, 1144051200, 1144054800, 1144058400, 
    1144062000, 1144065600, 1144069200, 1144072800, 1144076400, 1144080000, 
    1144083600, 1144087200, 1144090800, 1144094400, 1144098000, 1144101600, 
    1144105200, 1144108800, 1144112400, 1144116000, 1144119600, 1144123200, 
    1144126800, 1144130400, 1144134000, 1144137600, 1144141200, 1144144800, 
    1144148400, 1144152000, 1144155600, 1144159200, 1144162800, 1144166400, 
    1144170000, 1144173600, 1144177200, 1144180800, 1144184400, 1144188000, 
    1144191600, 1144195200, 1144198800, 1144202400, 1144206000, 1144209600, 
    1144213200, 1144216800, 1144220400, 1144224000, 1144227600, 1144231200, 
    1144234800, 1144238400, 1144242000, 1144245600, 1144249200, 1144252800, 
    1144256400, 1144260000, 1144263600, 1144267200, 1144270800, 1144274400, 
    1144278000, 1144281600, 1144285200, 1144288800, 1144292400, 1144296000, 
    1144299600, 1144303200, 1144306800, 1144310400, 1144314000, 1144317600, 
    1144321200, 1144324800, 1144328400, 1144332000, 1144335600, 1144339200, 
    1144342800, 1144346400, 1144350000, 1144353600, 1144357200, 1144360800, 
    1144364400, 1144368000, 1144371600, 1144375200, 1144378800, 1144382400, 
    1144386000, 1144389600, 1144393200, 1144396800, 1144400400, 1144404000, 
    1144407600, 1144411200, 1144414800, 1144418400, 1144422000, 1144425600, 
    1144429200, 1144432800, 1144436400, 1144440000, 1144443600, 1144447200, 
    1144450800, 1144454400, 1144458000, 1144461600, 1144465200, 1144468800, 
    1144472400, 1144476000, 1144479600, 1144483200, 1144486800, 1144490400, 
    1144494000, 1144497600, 1144501200, 1144504800, 1144508400, 1144512000, 
    1144515600, 1144519200, 1144522800, 1144526400, 1144530000, 1144533600, 
    1144537200, 1144540800, 1144544400, 1144548000, 1144551600, 1144555200, 
    1144558800, 1144562400, 1144566000, 1144569600, 1144573200, 1144576800, 
    1144580400, 1144584000, 1144587600, 1144591200, 1144594800, 1144598400, 
    1144602000, 1144605600, 1144609200, 1144612800, 1144616400, 1144620000, 
    1144623600, 1144627200, 1144630800, 1144634400, 1144638000, 1144641600, 
    1144645200, 1144648800, 1144652400, 1144656000, 1144659600, 1144663200, 
    1144666800, 1144670400, 1144674000, 1144677600, 1144681200, 1144684800, 
    1144688400, 1144692000, 1144695600, 1144699200, 1144702800, 1144706400, 
    1144710000, 1144713600, 1144717200, 1144720800, 1144724400, 1144728000, 
    1144731600, 1144735200, 1144738800, 1144742400, 1144746000, 1144749600, 
    1144753200, 1144756800, 1144760400, 1144764000, 1144767600, 1144771200, 
    1144774800, 1144778400, 1144782000, 1144785600, 1144789200, 1144792800, 
    1144796400, 1144800000, 1144803600, 1144807200, 1144810800, 1144814400, 
    1144818000, 1144821600, 1144825200, 1144828800, 1144832400, 1144836000, 
    1144839600, 1144843200, 1144846800, 1144850400, 1144854000, 1144857600, 
    1144861200, 1144864800, 1144868400, 1144872000, 1144875600, 1144879200, 
    1144882800, 1144886400, 1144890000, 1144893600, 1144897200, 1144900800, 
    1144904400, 1144908000, 1144911600, 1144915200, 1144918800, 1144922400, 
    1144926000, 1144929600, 1144933200, 1144936800, 1144940400, 1144944000, 
    1144947600, 1144951200, 1144954800, 1144958400, 1144962000, 1144965600, 
    1144969200, 1144972800, 1144976400, 1144980000, 1144983600, 1144987200, 
    1144990800, 1144994400, 1144998000, 1145001600, 1145005200, 1145008800, 
    1145012400, 1145016000, 1145019600, 1145023200, 1145026800, 1145030400, 
    1145034000, 1145037600, 1145041200, 1145044800, 1145048400, 1145052000, 
    1145055600, 1145059200, 1145062800, 1145066400, 1145070000, 1145073600, 
    1145077200, 1145080800, 1145084400, 1145088000, 1145091600, 1145095200, 
    1145098800, 1145102400, 1145106000, 1145109600, 1145113200, 1145116800, 
    1145120400, 1145124000, 1145127600, 1145131200, 1145134800, 1145138400, 
    1145142000, 1145145600, 1145149200, 1145152800, 1145156400, 1145160000, 
    1145163600, 1145167200, 1145170800, 1145174400, 1145178000, 1145181600, 
    1145185200, 1145188800, 1145192400, 1145196000, 1145199600, 1145203200, 
    1145206800, 1145210400, 1145214000, 1145217600, 1145221200, 1145224800, 
    1145228400, 1145232000, 1145235600, 1145239200, 1145242800, 1145246400, 
    1145250000, 1145253600, 1145257200, 1145260800, 1145264400, 1145268000, 
    1145271600, 1145275200, 1145278800, 1145282400, 1145286000, 1145289600, 
    1145293200, 1145296800, 1145300400, 1145304000, 1145307600, 1145311200, 
    1145314800, 1145318400, 1145322000, 1145325600, 1145329200, 1145332800, 
    1145336400, 1145340000, 1145343600, 1145347200, 1145350800, 1145354400, 
    1145358000, 1145361600, 1145365200, 1145368800, 1145372400, 1145376000, 
    1145379600, 1145383200, 1145386800, 1145390400, 1145394000, 1145397600, 
    1145401200, 1145404800, 1145408400, 1145412000, 1145415600, 1145419200, 
    1145422800, 1145426400, 1145430000, 1145433600, 1145437200, 1145440800, 
    1145444400, 1145448000, 1145451600, 1145455200, 1145458800, 1145462400, 
    1145466000, 1145469600, 1145473200, 1145476800, 1145480400, 1145484000, 
    1145487600, 1145491200, 1145494800, 1145498400, 1145502000, 1145505600, 
    1145509200, 1145512800, 1145516400, 1145520000, 1145523600, 1145527200, 
    1145530800, 1145534400, 1145538000, 1145541600, 1145545200, 1145548800, 
    1145552400, 1145556000, 1145559600, 1145563200, 1145566800, 1145570400, 
    1145574000, 1145577600, 1145581200, 1145584800, 1145588400, 1145592000, 
    1145595600, 1145599200, 1145602800, 1145606400, 1145610000, 1145613600, 
    1145617200, 1145620800, 1145624400, 1145628000, 1145631600, 1145635200, 
    1145638800, 1145642400, 1145646000, 1145649600, 1145653200, 1145656800, 
    1145660400, 1145664000, 1145667600, 1145671200, 1145674800, 1145678400, 
    1145682000, 1145685600, 1145689200, 1145692800, 1145696400, 1145700000, 
    1145703600, 1145707200, 1145710800, 1145714400, 1145718000, 1145721600, 
    1145725200, 1145728800, 1145732400, 1145736000, 1145739600, 1145743200, 
    1145746800, 1145750400, 1145754000, 1145757600, 1145761200, 1145764800, 
    1145768400, 1145772000, 1145775600, 1145779200, 1145782800, 1145786400, 
    1145790000, 1145793600, 1145797200, 1145800800, 1145804400, 1145808000, 
    1145811600, 1145815200, 1145818800, 1145822400, 1145826000, 1145829600, 
    1145833200, 1145836800, 1145840400, 1145844000, 1145847600, 1145851200, 
    1145854800, 1145858400, 1145862000, 1145865600, 1145869200, 1145872800, 
    1145876400, 1145880000, 1145883600, 1145887200, 1145890800, 1145894400, 
    1145898000, 1145901600, 1145905200, 1145908800, 1145912400, 1145916000, 
    1145919600, 1145923200, 1145926800, 1145930400, 1145934000, 1145937600, 
    1145941200, 1145944800, 1145948400, 1145952000, 1145955600, 1145959200, 
    1145962800, 1145966400, 1145970000, 1145973600, 1145977200, 1145980800, 
    1145984400, 1145988000, 1145991600, 1145995200, 1145998800, 1146002400, 
    1146006000, 1146009600, 1146013200, 1146016800, 1146020400, 1146024000, 
    1146027600, 1146031200, 1146034800, 1146038400, 1146042000, 1146045600, 
    1146049200, 1146052800, 1146056400, 1146060000, 1146063600, 1146067200, 
    1146070800, 1146074400, 1146078000, 1146081600, 1146085200, 1146088800, 
    1146092400, 1146096000, 1146099600, 1146103200, 1146106800, 1146110400, 
    1146114000, 1146117600, 1146121200, 1146124800, 1146128400, 1146132000, 
    1146135600, 1146139200, 1146142800, 1146146400, 1146150000, 1146153600, 
    1146157200, 1146160800, 1146164400, 1146168000, 1146171600, 1146175200, 
    1146178800, 1146182400, 1146186000, 1146189600, 1146193200, 1146196800, 
    1146200400, 1146204000, 1146207600, 1146211200, 1146214800, 1146218400, 
    1146222000, 1146225600, 1146229200, 1146232800, 1146236400, 1146240000, 
    1146243600, 1146247200, 1146250800, 1146254400, 1146258000, 1146261600, 
    1146265200, 1146268800, 1146272400, 1146276000, 1146279600, 1146283200, 
    1146286800, 1146290400, 1146294000, 1146297600, 1146301200, 1146304800, 
    1146308400, 1146312000, 1146315600, 1146319200, 1146322800, 1146326400, 
    1146330000, 1146333600, 1146337200, 1146340800, 1146344400, 1146348000, 
    1146351600, 1146355200, 1146358800, 1146362400, 1146366000, 1146369600, 
    1146373200, 1146376800, 1146380400, 1146384000, 1146387600, 1146391200, 
    1146394800, 1146398400, 1146402000, 1146405600, 1146409200, 1146412800, 
    1146416400, 1146420000, 1146423600, 1146427200, 1146430800, 1146434400, 
    1146438000, 1146441600, 1146445200, 1146448800, 1146452400, 1146456000, 
    1146459600, 1146463200, 1146466800, 1146470400, 1146474000, 1146477600, 
    1146481200, 1146484800, 1146488400, 1146492000, 1146495600, 1146499200, 
    1146502800, 1146506400, 1146510000, 1146513600, 1146517200, 1146520800, 
    1146524400, 1146528000, 1146531600, 1146535200, 1146538800, 1146542400, 
    1146546000, 1146549600, 1146553200, 1146556800, 1146560400, 1146564000, 
    1146567600, 1146571200, 1146574800, 1146578400, 1146582000, 1146585600, 
    1146589200, 1146592800, 1146596400, 1146600000, 1146603600, 1146607200, 
    1146610800, 1146614400, 1146618000, 1146621600, 1146625200, 1146628800, 
    1146632400, 1146636000, 1146639600, 1146643200, 1146646800, 1146650400, 
    1146654000, 1146657600, 1146661200, 1146664800, 1146668400, 1146672000, 
    1146675600, 1146679200, 1146682800, 1146686400, 1146690000, 1146693600, 
    1146697200, 1146700800, 1146704400, 1146708000, 1146711600, 1146715200, 
    1146718800, 1146722400, 1146726000, 1146729600, 1146733200, 1146736800, 
    1146740400, 1146744000, 1146747600, 1146751200, 1146754800, 1146758400, 
    1146762000, 1146765600, 1146769200, 1146772800, 1146776400, 1146780000, 
    1146783600, 1146787200, 1146790800, 1146794400, 1146798000, 1146801600, 
    1146805200, 1146808800, 1146812400, 1146816000, 1146819600, 1146823200, 
    1146826800, 1146830400, 1146834000, 1146837600, 1146841200, 1146844800, 
    1146848400, 1146852000, 1146855600, 1146859200, 1146862800, 1146866400, 
    1146870000, 1146873600, 1146877200, 1146880800, 1146884400, 1146888000, 
    1146891600, 1146895200, 1146898800, 1146902400, 1146906000, 1146909600, 
    1146913200, 1146916800, 1146920400, 1146924000, 1146927600, 1146931200, 
    1146934800, 1146938400, 1146942000, 1146945600, 1146949200, 1146952800, 
    1146956400, 1146960000, 1146963600, 1146967200, 1146970800, 1146974400, 
    1146978000, 1146981600, 1146985200, 1146988800, 1146992400, 1146996000, 
    1146999600, 1147003200, 1147006800, 1147010400, 1147014000, 1147017600, 
    1147021200, 1147024800, 1147028400, 1147032000, 1147035600, 1147039200, 
    1147042800, 1147046400, 1147050000, 1147053600, 1147057200, 1147060800, 
    1147064400, 1147068000, 1147071600, 1147075200, 1147078800, 1147082400, 
    1147086000, 1147089600, 1147093200, 1147096800, 1147100400, 1147104000, 
    1147107600, 1147111200, 1147114800, 1147118400, 1147122000, 1147125600, 
    1147129200, 1147132800, 1147136400, 1147140000, 1147143600, 1147147200, 
    1147150800, 1147154400, 1147158000, 1147161600, 1147165200, 1147168800, 
    1147172400, 1147176000, 1147179600, 1147183200, 1147186800, 1147190400, 
    1147194000, 1147197600, 1147201200, 1147204800, 1147208400, 1147212000, 
    1147215600, 1147219200, 1147222800, 1147226400, 1147230000, 1147233600, 
    1147237200, 1147240800, 1147244400, 1147248000, 1147251600, 1147255200, 
    1147258800, 1147262400, 1147266000, 1147269600, 1147273200, 1147276800, 
    1147280400, 1147284000, 1147287600, 1147291200, 1147294800, 1147298400, 
    1147302000, 1147305600, 1147309200, 1147312800, 1147316400, 1147320000, 
    1147323600, 1147327200, 1147330800, 1147334400, 1147338000, 1147341600, 
    1147345200, 1147348800, 1147352400, 1147356000, 1147359600, 1147363200, 
    1147366800, 1147370400, 1147374000, 1147377600, 1147381200, 1147384800, 
    1147388400, 1147392000, 1147395600, 1147399200, 1147402800, 1147406400, 
    1147410000, 1147413600, 1147417200, 1147420800, 1147424400, 1147428000, 
    1147431600, 1147435200, 1147438800, 1147442400, 1147446000, 1147449600, 
    1147453200, 1147456800, 1147460400, 1147464000, 1147467600, 1147471200, 
    1147474800, 1147478400, 1147482000, 1147485600, 1147489200, 1147492800, 
    1147496400, 1147500000, 1147503600, 1147507200, 1147510800, 1147514400, 
    1147518000, 1147521600, 1147525200, 1147528800, 1147532400, 1147536000, 
    1147539600, 1147543200, 1147546800, 1147550400, 1147554000, 1147557600, 
    1147561200, 1147564800, 1147568400, 1147572000, 1147575600, 1147579200, 
    1147582800, 1147586400, 1147590000, 1147593600, 1147597200, 1147600800, 
    1147604400, 1147608000, 1147611600, 1147615200, 1147618800, 1147622400, 
    1147626000, 1147629600, 1147633200, 1147636800, 1147640400, 1147644000, 
    1147647600, 1147651200, 1147654800, 1147658400, 1147662000, 1147665600, 
    1147669200, 1147672800, 1147676400, 1147680000, 1147683600, 1147687200, 
    1147690800, 1147694400, 1147698000, 1147701600, 1147705200, 1147708800, 
    1147712400, 1147716000, 1147719600, 1147723200, 1147726800, 1147730400, 
    1147734000, 1147737600, 1147741200, 1147744800, 1147748400, 1147752000, 
    1147755600, 1147759200, 1147762800, 1147766400, 1147770000, 1147773600, 
    1147777200, 1147780800, 1147784400, 1147788000, 1147791600, 1147795200, 
    1147798800, 1147802400, 1147806000, 1147809600, 1147813200, 1147816800, 
    1147820400, 1147824000, 1147827600, 1147831200, 1147834800, 1147838400, 
    1147842000, 1147845600, 1147849200, 1147852800, 1147856400, 1147860000, 
    1147863600, 1147867200, 1147870800, 1147874400, 1147878000, 1147881600, 
    1147885200, 1147888800, 1147892400, 1147896000, 1147899600, 1147903200, 
    1147906800, 1147910400, 1147914000, 1147917600, 1147921200, 1147924800, 
    1147928400, 1147932000, 1147935600, 1147939200, 1147942800, 1147946400, 
    1147950000, 1147953600, 1147957200, 1147960800, 1147964400, 1147968000, 
    1147971600, 1147975200, 1147978800, 1147982400, 1147986000, 1147989600, 
    1147993200, 1147996800, 1148000400, 1148004000, 1148007600, 1148011200, 
    1148014800, 1148018400, 1148022000, 1148025600, 1148029200, 1148032800, 
    1148036400, 1148040000, 1148043600, 1148047200, 1148050800, 1148054400, 
    1148058000, 1148061600, 1148065200, 1148068800, 1148072400, 1148076000, 
    1148079600, 1148083200, 1148086800, 1148090400, 1148094000, 1148097600, 
    1148101200, 1148104800, 1148108400, 1148112000, 1148115600, 1148119200, 
    1148122800, 1148126400, 1148130000, 1148133600, 1148137200, 1148140800, 
    1148144400, 1148148000, 1148151600, 1148155200, 1148158800, 1148162400, 
    1148166000, 1148169600, 1148173200, 1148176800, 1148180400, 1148184000, 
    1148187600, 1148191200, 1148194800, 1148198400, 1148202000, 1148205600, 
    1148209200, 1148212800, 1148216400, 1148220000, 1148223600, 1148227200, 
    1148230800, 1148234400, 1148238000, 1148241600, 1148245200, 1148248800, 
    1148252400, 1148256000, 1148259600, 1148263200, 1148266800, 1148270400, 
    1148274000, 1148277600, 1148281200, 1148284800, 1148288400, 1148292000, 
    1148295600, 1148299200, 1148302800, 1148306400, 1148310000, 1148313600, 
    1148317200, 1148320800, 1148324400, 1148328000, 1148331600, 1148335200, 
    1148338800, 1148342400, 1148346000, 1148349600, 1148353200, 1148356800, 
    1148360400, 1148364000, 1148367600, 1148371200, 1148374800, 1148378400, 
    1148382000, 1148385600, 1148389200, 1148392800, 1148396400, 1148400000, 
    1148403600, 1148407200, 1148410800, 1148414400, 1148418000, 1148421600, 
    1148425200, 1148428800, 1148432400, 1148436000, 1148439600, 1148443200, 
    1148446800, 1148450400, 1148454000, 1148457600, 1148461200, 1148464800, 
    1148468400, 1148472000, 1148475600, 1148479200, 1148482800, 1148486400, 
    1148490000, 1148493600, 1148497200, 1148500800, 1148504400, 1148508000, 
    1148511600, 1148515200, 1148518800, 1148522400, 1148526000, 1148529600, 
    1148533200, 1148536800, 1148540400, 1148544000, 1148547600, 1148551200, 
    1148554800, 1148558400, 1148562000, 1148565600, 1148569200, 1148572800, 
    1148576400, 1148580000, 1148583600, 1148587200, 1148590800, 1148594400, 
    1148598000, 1148601600, 1148605200, 1148608800, 1148612400, 1148616000, 
    1148619600, 1148623200, 1148626800, 1148630400, 1148634000, 1148637600, 
    1148641200, 1148644800, 1148648400, 1148652000, 1148655600, 1148659200, 
    1148662800, 1148666400, 1148670000, 1148673600, 1148677200, 1148680800, 
    1148684400, 1148688000, 1148691600, 1148695200, 1148698800, 1148702400, 
    1148706000, 1148709600, 1148713200, 1148716800, 1148720400, 1148724000, 
    1148727600, 1148731200, 1148734800, 1148738400, 1148742000, 1148745600, 
    1148749200, 1148752800, 1148756400, 1148760000, 1148763600, 1148767200, 
    1148770800, 1148774400, 1148778000, 1148781600, 1148785200, 1148788800, 
    1148792400, 1148796000, 1148799600, 1148803200, 1148806800, 1148810400, 
    1148814000, 1148817600, 1148821200, 1148824800, 1148828400, 1148832000, 
    1148835600, 1148839200, 1148842800, 1148846400, 1148850000, 1148853600, 
    1148857200, 1148860800, 1148864400, 1148868000, 1148871600, 1148875200, 
    1148878800, 1148882400, 1148886000, 1148889600, 1148893200, 1148896800, 
    1148900400, 1148904000, 1148907600, 1148911200, 1148914800, 1148918400, 
    1148922000, 1148925600, 1148929200, 1148932800, 1148936400, 1148940000, 
    1148943600, 1148947200, 1148950800, 1148954400, 1148958000, 1148961600, 
    1148965200, 1148968800, 1148972400, 1148976000, 1148979600, 1148983200, 
    1148986800, 1148990400, 1148994000, 1148997600, 1149001200, 1149004800, 
    1149008400, 1149012000, 1149015600, 1149019200, 1149022800, 1149026400, 
    1149030000, 1149033600, 1149037200, 1149040800, 1149044400, 1149048000, 
    1149051600, 1149055200, 1149058800, 1149062400, 1149066000, 1149069600, 
    1149073200, 1149076800, 1149080400, 1149084000, 1149087600, 1149091200, 
    1149094800, 1149098400, 1149102000, 1149105600, 1149109200, 1149112800, 
    1149116400, 1149120000, 1149123600, 1149127200, 1149130800, 1149134400, 
    1149138000, 1149141600, 1149145200, 1149148800, 1149152400, 1149156000, 
    1149159600, 1149163200, 1149166800, 1149170400, 1149174000, 1149177600, 
    1149181200, 1149184800, 1149188400, 1149192000, 1149195600, 1149199200, 
    1149202800, 1149206400, 1149210000, 1149213600, 1149217200, 1149220800, 
    1149224400, 1149228000, 1149231600, 1149235200, 1149238800, 1149242400, 
    1149246000, 1149249600, 1149253200, 1149256800, 1149260400, 1149264000, 
    1149267600, 1149271200, 1149274800, 1149278400, 1149282000, 1149285600, 
    1149289200, 1149292800, 1149296400, 1149300000, 1149303600, 1149307200, 
    1149310800, 1149314400, 1149318000, 1149321600, 1149325200, 1149328800, 
    1149332400, 1149336000, 1149339600, 1149343200, 1149346800, 1149350400, 
    1149354000, 1149357600, 1149361200, 1149364800, 1149368400, 1149372000, 
    1149375600, 1149379200, 1149382800, 1149386400, 1149390000, 1149393600, 
    1149397200, 1149400800, 1149404400, 1149408000, 1149411600, 1149415200, 
    1149418800, 1149422400, 1149426000, 1149429600, 1149433200, 1149436800, 
    1149440400, 1149444000, 1149447600, 1149451200, 1149454800, 1149458400, 
    1149462000, 1149465600, 1149469200, 1149472800, 1149476400, 1149480000, 
    1149483600, 1149487200, 1149490800, 1149494400, 1149498000, 1149501600, 
    1149505200, 1149508800, 1149512400, 1149516000, 1149519600, 1149523200, 
    1149526800, 1149530400, 1149534000, 1149537600, 1149541200, 1149544800, 
    1149548400, 1149552000, 1149555600, 1149559200, 1149562800, 1149566400, 
    1149570000, 1149573600, 1149577200, 1149580800, 1149584400, 1149588000, 
    1149591600, 1149595200, 1149598800, 1149602400, 1149606000, 1149609600, 
    1149613200, 1149616800, 1149620400, 1149624000, 1149627600, 1149631200, 
    1149634800, 1149638400, 1149642000, 1149645600, 1149649200, 1149652800, 
    1149656400, 1149660000, 1149663600, 1149667200, 1149670800, 1149674400, 
    1149678000, 1149681600, 1149685200, 1149688800, 1149692400, 1149696000, 
    1149699600, 1149703200, 1149706800, 1149710400, 1149714000, 1149717600, 
    1149721200, 1149724800, 1149728400, 1149732000, 1149735600, 1149739200, 
    1149742800, 1149746400, 1149750000, 1149753600, 1149757200, 1149760800, 
    1149764400, 1149768000, 1149771600, 1149775200, 1149778800, 1149782400, 
    1149786000, 1149789600, 1149793200, 1149796800, 1149800400, 1149804000, 
    1149807600, 1149811200, 1149814800, 1149818400, 1149822000, 1149825600, 
    1149829200, 1149832800, 1149836400, 1149840000, 1149843600, 1149847200, 
    1149850800, 1149854400, 1149858000, 1149861600, 1149865200, 1149868800, 
    1149872400, 1149876000, 1149879600, 1149883200, 1149886800, 1149890400, 
    1149894000, 1149897600, 1149901200, 1149904800, 1149908400, 1149912000, 
    1149915600, 1149919200, 1149922800, 1149926400, 1149930000, 1149933600, 
    1149937200, 1149940800, 1149944400, 1149948000, 1149951600, 1149955200, 
    1149958800, 1149962400, 1149966000, 1149969600, 1149973200, 1149976800, 
    1149980400, 1149984000, 1149987600, 1149991200, 1149994800, 1149998400, 
    1150002000, 1150005600, 1150009200, 1150012800, 1150016400, 1150020000, 
    1150023600, 1150027200, 1150030800, 1150034400, 1150038000, 1150041600, 
    1150045200, 1150048800, 1150052400, 1150056000, 1150059600, 1150063200, 
    1150066800, 1150070400, 1150074000, 1150077600, 1150081200, 1150084800, 
    1150088400, 1150092000, 1150095600, 1150099200, 1150102800, 1150106400, 
    1150110000, 1150113600, 1150117200, 1150120800, 1150124400, 1150128000, 
    1150131600, 1150135200, 1150138800, 1150142400, 1150146000, 1150149600, 
    1150153200, 1150156800, 1150160400, 1150164000, 1150167600, 1150171200, 
    1150174800, 1150178400, 1150182000, 1150185600, 1150189200, 1150192800, 
    1150196400, 1150200000, 1150203600, 1150207200, 1150210800, 1150214400, 
    1150218000, 1150221600, 1150225200, 1150228800, 1150232400, 1150236000, 
    1150239600, 1150243200, 1150246800, 1150250400, 1150254000, 1150257600, 
    1150261200, 1150264800, 1150268400, 1150272000, 1150275600, 1150279200, 
    1150282800, 1150286400, 1150290000, 1150293600, 1150297200, 1150300800, 
    1150304400, 1150308000, 1150311600, 1150315200, 1150318800, 1150322400, 
    1150326000, 1150329600, 1150333200, 1150336800, 1150340400, 1150344000, 
    1150347600, 1150351200, 1150354800, 1150358400, 1150362000, 1150365600, 
    1150369200, 1150372800, 1150376400, 1150380000, 1150383600, 1150387200, 
    1150390800, 1150394400, 1150398000, 1150401600, 1150405200, 1150408800, 
    1150412400, 1150416000, 1150419600, 1150423200, 1150426800, 1150430400, 
    1150434000, 1150437600, 1150441200, 1150444800, 1150448400, 1150452000, 
    1150455600, 1150459200, 1150462800, 1150466400, 1150470000, 1150473600, 
    1150477200, 1150480800, 1150484400, 1150488000, 1150491600, 1150495200, 
    1150498800, 1150502400, 1150506000, 1150509600, 1150513200, 1150516800, 
    1150520400, 1150524000, 1150527600, 1150531200, 1150534800, 1150538400, 
    1150542000, 1150545600, 1150549200, 1150552800, 1150556400, 1150560000, 
    1150563600, 1150567200, 1150570800, 1150574400, 1150578000, 1150581600, 
    1150585200, 1150588800, 1150592400, 1150596000, 1150599600, 1150603200, 
    1150606800, 1150610400, 1150614000, 1150617600, 1150621200, 1150624800, 
    1150628400, 1150632000, 1150635600, 1150639200, 1150642800, 1150646400, 
    1150650000, 1150653600, 1150657200, 1150660800, 1150664400, 1150668000, 
    1150671600, 1150675200, 1150678800, 1150682400, 1150686000, 1150689600, 
    1150693200, 1150696800, 1150700400, 1150704000, 1150707600, 1150711200, 
    1150714800, 1150718400, 1150722000, 1150725600, 1150729200, 1150732800, 
    1150736400, 1150740000, 1150743600, 1150747200, 1150750800, 1150754400, 
    1150758000, 1150761600, 1150765200, 1150768800, 1150772400, 1150776000, 
    1150779600, 1150783200, 1150786800, 1150790400, 1150794000, 1150797600, 
    1150801200, 1150804800, 1150808400, 1150812000, 1150815600, 1150819200, 
    1150822800, 1150826400, 1150830000, 1150833600, 1150837200, 1150840800, 
    1150844400, 1150848000, 1150851600, 1150855200, 1150858800, 1150862400, 
    1150866000, 1150869600, 1150873200, 1150876800, 1150880400, 1150884000, 
    1150887600, 1150891200, 1150894800, 1150898400, 1150902000, 1150905600, 
    1150909200, 1150912800, 1150916400, 1150920000, 1150923600, 1150927200, 
    1150930800, 1150934400, 1150938000, 1150941600, 1150945200, 1150948800, 
    1150952400, 1150956000, 1150959600, 1150963200, 1150966800, 1150970400, 
    1150974000, 1150977600, 1150981200, 1150984800, 1150988400, 1150992000, 
    1150995600, 1150999200, 1151002800, 1151006400, 1151010000, 1151013600, 
    1151017200, 1151020800, 1151024400, 1151028000, 1151031600, 1151035200, 
    1151038800, 1151042400, 1151046000, 1151049600, 1151053200, 1151056800, 
    1151060400, 1151064000, 1151067600, 1151071200, 1151074800, 1151078400, 
    1151082000, 1151085600, 1151089200, 1151092800, 1151096400, 1151100000, 
    1151103600, 1151107200, 1151110800, 1151114400, 1151118000, 1151121600, 
    1151125200, 1151128800, 1151132400, 1151136000, 1151139600, 1151143200, 
    1151146800, 1151150400, 1151154000, 1151157600, 1151161200, 1151164800, 
    1151168400, 1151172000, 1151175600, 1151179200, 1151182800, 1151186400, 
    1151190000, 1151193600, 1151197200, 1151200800, 1151204400, 1151208000, 
    1151211600, 1151215200, 1151218800, 1151222400, 1151226000, 1151229600, 
    1151233200, 1151236800, 1151240400, 1151244000, 1151247600, 1151251200, 
    1151254800, 1151258400, 1151262000, 1151265600, 1151269200, 1151272800, 
    1151276400, 1151280000, 1151283600, 1151287200, 1151290800, 1151294400, 
    1151298000, 1151301600, 1151305200, 1151308800, 1151312400, 1151316000, 
    1151319600, 1151323200, 1151326800, 1151330400, 1151334000, 1151337600, 
    1151341200, 1151344800, 1151348400, 1151352000, 1151355600, 1151359200, 
    1151362800, 1151366400, 1151370000, 1151373600, 1151377200, 1151380800, 
    1151384400, 1151388000, 1151391600, 1151395200, 1151398800, 1151402400, 
    1151406000, 1151409600, 1151413200, 1151416800, 1151420400, 1151424000, 
    1151427600, 1151431200, 1151434800, 1151438400, 1151442000, 1151445600, 
    1151449200, 1151452800, 1151456400, 1151460000, 1151463600, 1151467200, 
    1151470800, 1151474400, 1151478000, 1151481600, 1151485200, 1151488800, 
    1151492400, 1151496000, 1151499600, 1151503200, 1151506800, 1151510400, 
    1151514000, 1151517600, 1151521200, 1151524800, 1151528400, 1151532000, 
    1151535600, 1151539200, 1151542800, 1151546400, 1151550000, 1151553600, 
    1151557200, 1151560800, 1151564400, 1151568000, 1151571600, 1151575200, 
    1151578800, 1151582400, 1151586000, 1151589600, 1151593200, 1151596800, 
    1151600400, 1151604000, 1151607600, 1151611200, 1151614800, 1151618400, 
    1151622000, 1151625600, 1151629200, 1151632800, 1151636400, 1151640000, 
    1151643600, 1151647200, 1151650800, 1151654400, 1151658000, 1151661600, 
    1151665200, 1151668800, 1151672400, 1151676000, 1151679600, 1151683200, 
    1151686800, 1151690400, 1151694000, 1151697600, 1151701200, 1151704800, 
    1151708400, 1151712000, 1151715600, 1151719200, 1151722800, 1151726400, 
    1151730000, 1151733600, 1151737200, 1151740800, 1151744400, 1151748000, 
    1151751600, 1151755200, 1151758800, 1151762400, 1151766000, 1151769600, 
    1151773200, 1151776800, 1151780400, 1151784000, 1151787600, 1151791200, 
    1151794800, 1151798400, 1151802000, 1151805600, 1151809200, 1151812800, 
    1151816400, 1151820000, 1151823600, 1151827200, 1151830800, 1151834400, 
    1151838000, 1151841600, 1151845200, 1151848800, 1151852400, 1151856000, 
    1151859600, 1151863200, 1151866800, 1151870400, 1151874000, 1151877600, 
    1151881200, 1151884800, 1151888400, 1151892000, 1151895600, 1151899200, 
    1151902800, 1151906400, 1151910000, 1151913600, 1151917200, 1151920800, 
    1151924400, 1151928000, 1151931600, 1151935200, 1151938800, 1151942400, 
    1151946000, 1151949600, 1151953200, 1151956800, 1151960400, 1151964000, 
    1151967600, 1151971200, 1151974800, 1151978400, 1151982000, 1151985600, 
    1151989200, 1151992800, 1151996400, 1152000000, 1152003600, 1152007200, 
    1152010800, 1152014400, 1152018000, 1152021600, 1152025200, 1152028800, 
    1152032400, 1152036000, 1152039600, 1152043200, 1152046800, 1152050400, 
    1152054000, 1152057600, 1152061200, 1152064800, 1152068400, 1152072000, 
    1152075600, 1152079200, 1152082800, 1152086400, 1152090000, 1152093600, 
    1152097200, 1152100800, 1152104400, 1152108000, 1152111600, 1152115200, 
    1152118800, 1152122400, 1152126000, 1152129600, 1152133200, 1152136800, 
    1152140400, 1152144000, 1152147600, 1152151200, 1152154800, 1152158400, 
    1152162000, 1152165600, 1152169200, 1152172800, 1152176400, 1152180000, 
    1152183600, 1152187200, 1152190800, 1152194400, 1152198000, 1152201600, 
    1152205200, 1152208800, 1152212400, 1152216000, 1152219600, 1152223200, 
    1152226800, 1152230400, 1152234000, 1152237600, 1152241200, 1152244800, 
    1152248400, 1152252000, 1152255600, 1152259200, 1152262800, 1152266400, 
    1152270000, 1152273600, 1152277200, 1152280800, 1152284400, 1152288000, 
    1152291600, 1152295200, 1152298800, 1152302400, 1152306000, 1152309600, 
    1152313200, 1152316800, 1152320400, 1152324000, 1152327600, 1152331200, 
    1152334800, 1152338400, 1152342000, 1152345600, 1152349200, 1152352800, 
    1152356400, 1152360000, 1152363600, 1152367200, 1152370800, 1152374400, 
    1152378000, 1152381600, 1152385200, 1152388800, 1152392400, 1152396000, 
    1152399600, 1152403200, 1152406800, 1152410400, 1152414000, 1152417600, 
    1152421200, 1152424800, 1152428400, 1152432000, 1152435600, 1152439200, 
    1152442800, 1152446400, 1152450000, 1152453600, 1152457200, 1152460800, 
    1152464400, 1152468000, 1152471600, 1152475200, 1152478800, 1152482400, 
    1152486000, 1152489600, 1152493200, 1152496800, 1152500400, 1152504000, 
    1152507600, 1152511200, 1152514800, 1152518400, 1152522000, 1152525600, 
    1152529200, 1152532800, 1152536400, 1152540000, 1152543600, 1152547200, 
    1152550800, 1152554400, 1152558000, 1152561600, 1152565200, 1152568800, 
    1152572400, 1152576000, 1152579600, 1152583200, 1152586800, 1152590400, 
    1152594000, 1152597600, 1152601200, 1152604800, 1152608400, 1152612000, 
    1152615600, 1152619200, 1152622800, 1152626400, 1152630000, 1152633600, 
    1152637200, 1152640800, 1152644400, 1152648000, 1152651600, 1152655200, 
    1152658800, 1152662400, 1152666000, 1152669600, 1152673200, 1152676800, 
    1152680400, 1152684000, 1152687600, 1152691200, 1152694800, 1152698400, 
    1152702000, 1152705600, 1152709200, 1152712800, 1152716400, 1152720000, 
    1152723600, 1152727200, 1152730800, 1152734400, 1152738000, 1152741600, 
    1152745200, 1152748800, 1152752400, 1152756000, 1152759600, 1152763200, 
    1152766800, 1152770400, 1152774000, 1152777600, 1152781200, 1152784800, 
    1152788400, 1152792000, 1152795600, 1152799200, 1152802800, 1152806400, 
    1152810000, 1152813600, 1152817200, 1152820800, 1152824400, 1152828000, 
    1152831600, 1152835200, 1152838800, 1152842400, 1152846000, 1152849600, 
    1152853200, 1152856800, 1152860400, 1152864000, 1152867600, 1152871200, 
    1152874800, 1152878400, 1152882000, 1152885600, 1152889200, 1152892800, 
    1152896400, 1152900000, 1152903600, 1152907200, 1152910800, 1152914400, 
    1152918000, 1152921600, 1152925200, 1152928800, 1152932400, 1152936000, 
    1152939600, 1152943200, 1152946800, 1152950400, 1152954000, 1152957600, 
    1152961200, 1152964800, 1152968400, 1152972000, 1152975600, 1152979200, 
    1152982800, 1152986400, 1152990000, 1152993600, 1152997200, 1153000800, 
    1153004400, 1153008000, 1153011600, 1153015200, 1153018800, 1153022400, 
    1153026000, 1153029600, 1153033200, 1153036800, 1153040400, 1153044000, 
    1153047600, 1153051200, 1153054800, 1153058400, 1153062000, 1153065600, 
    1153069200, 1153072800, 1153076400, 1153080000, 1153083600, 1153087200, 
    1153090800, 1153094400, 1153098000, 1153101600, 1153105200, 1153108800, 
    1153112400, 1153116000, 1153119600, 1153123200, 1153126800, 1153130400, 
    1153134000, 1153137600, 1153141200, 1153144800, 1153148400, 1153152000, 
    1153155600, 1153159200, 1153162800, 1153166400, 1153170000, 1153173600, 
    1153177200, 1153180800, 1153184400, 1153188000, 1153191600, 1153195200, 
    1153198800, 1153202400, 1153206000, 1153209600, 1153213200, 1153216800, 
    1153220400, 1153224000, 1153227600, 1153231200, 1153234800, 1153238400, 
    1153242000, 1153245600, 1153249200, 1153252800, 1153256400, 1153260000, 
    1153263600, 1153267200, 1153270800, 1153274400, 1153278000, 1153281600, 
    1153285200, 1153288800, 1153292400, 1153296000, 1153299600, 1153303200, 
    1153306800, 1153310400, 1153314000, 1153317600, 1153321200, 1153324800, 
    1153328400, 1153332000, 1153335600, 1153339200, 1153342800, 1153346400, 
    1153350000, 1153353600, 1153357200, 1153360800, 1153364400, 1153368000, 
    1153371600, 1153375200, 1153378800, 1153382400, 1153386000, 1153389600, 
    1153393200, 1153396800, 1153400400, 1153404000, 1153407600, 1153411200, 
    1153414800, 1153418400, 1153422000, 1153425600, 1153429200, 1153432800, 
    1153436400, 1153440000, 1153443600, 1153447200, 1153450800, 1153454400, 
    1153458000, 1153461600, 1153465200, 1153468800, 1153472400, 1153476000, 
    1153479600, 1153483200, 1153486800, 1153490400, 1153494000, 1153497600, 
    1153501200, 1153504800, 1153508400, 1153512000, 1153515600, 1153519200, 
    1153522800, 1153526400, 1153530000, 1153533600, 1153537200, 1153540800, 
    1153544400, 1153548000, 1153551600, 1153555200, 1153558800, 1153562400, 
    1153566000, 1153569600, 1153573200, 1153576800, 1153580400, 1153584000, 
    1153587600, 1153591200, 1153594800, 1153598400, 1153602000, 1153605600, 
    1153609200, 1153612800, 1153616400, 1153620000, 1153623600, 1153627200, 
    1153630800, 1153634400, 1153638000, 1153641600, 1153645200, 1153648800, 
    1153652400, 1153656000, 1153659600, 1153663200, 1153666800, 1153670400, 
    1153674000, 1153677600, 1153681200, 1153684800, 1153688400, 1153692000, 
    1153695600, 1153699200, 1153702800, 1153706400, 1153710000, 1153713600, 
    1153717200, 1153720800, 1153724400, 1153728000, 1153731600, 1153735200, 
    1153738800, 1153742400, 1153746000, 1153749600, 1153753200, 1153756800, 
    1153760400, 1153764000, 1153767600, 1153771200, 1153774800, 1153778400, 
    1153782000, 1153785600, 1153789200, 1153792800, 1153796400, 1153800000, 
    1153803600, 1153807200, 1153810800, 1153814400, 1153818000, 1153821600, 
    1153825200, 1153828800, 1153832400, 1153836000, 1153839600, 1153843200, 
    1153846800, 1153850400, 1153854000, 1153857600, 1153861200, 1153864800, 
    1153868400, 1153872000, 1153875600, 1153879200, 1153882800, 1153886400, 
    1153890000, 1153893600, 1153897200, 1153900800, 1153904400, 1153908000, 
    1153911600, 1153915200, 1153918800, 1153922400, 1153926000, 1153929600, 
    1153933200, 1153936800, 1153940400, 1153944000, 1153947600, 1153951200, 
    1153954800, 1153958400, 1153962000, 1153965600, 1153969200, 1153972800, 
    1153976400, 1153980000, 1153983600, 1153987200, 1153990800, 1153994400, 
    1153998000, 1154001600, 1154005200, 1154008800, 1154012400, 1154016000, 
    1154019600, 1154023200, 1154026800, 1154030400, 1154034000, 1154037600, 
    1154041200, 1154044800, 1154048400, 1154052000, 1154055600, 1154059200, 
    1154062800, 1154066400, 1154070000, 1154073600, 1154077200, 1154080800, 
    1154084400, 1154088000, 1154091600, 1154095200, 1154098800, 1154102400, 
    1154106000, 1154109600, 1154113200, 1154116800, 1154120400, 1154124000, 
    1154127600, 1154131200, 1154134800, 1154138400, 1154142000, 1154145600, 
    1154149200, 1154152800, 1154156400, 1154160000, 1154163600, 1154167200, 
    1154170800, 1154174400, 1154178000, 1154181600, 1154185200, 1154188800, 
    1154192400, 1154196000, 1154199600, 1154203200, 1154206800, 1154210400, 
    1154214000, 1154217600, 1154221200, 1154224800, 1154228400, 1154232000, 
    1154235600, 1154239200, 1154242800, 1154246400, 1154250000, 1154253600, 
    1154257200, 1154260800, 1154264400, 1154268000, 1154271600, 1154275200, 
    1154278800, 1154282400, 1154286000, 1154289600, 1154293200, 1154296800, 
    1154300400, 1154304000, 1154307600, 1154311200, 1154314800, 1154318400, 
    1154322000, 1154325600, 1154329200, 1154332800, 1154336400, 1154340000, 
    1154343600, 1154347200, 1154350800, 1154354400, 1154358000, 1154361600, 
    1154365200, 1154368800, 1154372400, 1154376000, 1154379600, 1154383200, 
    1154386800, 1154390400, 1154394000, 1154397600, 1154401200, 1154404800, 
    1154408400, 1154412000, 1154415600, 1154419200, 1154422800, 1154426400, 
    1154430000, 1154433600, 1154437200, 1154440800, 1154444400, 1154448000, 
    1154451600, 1154455200, 1154458800, 1154462400, 1154466000, 1154469600, 
    1154473200, 1154476800, 1154480400, 1154484000, 1154487600, 1154491200, 
    1154494800, 1154498400, 1154502000, 1154505600, 1154509200, 1154512800, 
    1154516400, 1154520000, 1154523600, 1154527200, 1154530800, 1154534400, 
    1154538000, 1154541600, 1154545200, 1154548800, 1154552400, 1154556000, 
    1154559600, 1154563200, 1154566800, 1154570400, 1154574000, 1154577600, 
    1154581200, 1154584800, 1154588400, 1154592000, 1154595600, 1154599200, 
    1154602800, 1154606400, 1154610000, 1154613600, 1154617200, 1154620800, 
    1154624400, 1154628000, 1154631600, 1154635200, 1154638800, 1154642400, 
    1154646000, 1154649600, 1154653200, 1154656800, 1154660400, 1154664000, 
    1154667600, 1154671200, 1154674800, 1154678400, 1154682000, 1154685600, 
    1154689200, 1154692800, 1154696400, 1154700000, 1154703600, 1154707200, 
    1154710800, 1154714400, 1154718000, 1154721600, 1154725200, 1154728800, 
    1154732400, 1154736000, 1154739600, 1154743200, 1154746800, 1154750400, 
    1154754000, 1154757600, 1154761200, 1154764800, 1154768400, 1154772000, 
    1154775600, 1154779200, 1154782800, 1154786400, 1154790000, 1154793600, 
    1154797200, 1154800800, 1154804400, 1154808000, 1154811600, 1154815200, 
    1154818800, 1154822400, 1154826000, 1154829600, 1154833200, 1154836800, 
    1154840400, 1154844000, 1154847600, 1154851200, 1154854800, 1154858400, 
    1154862000, 1154865600, 1154869200, 1154872800, 1154876400, 1154880000, 
    1154883600, 1154887200, 1154890800, 1154894400, 1154898000, 1154901600, 
    1154905200, 1154908800, 1154912400, 1154916000, 1154919600, 1154923200, 
    1154926800, 1154930400, 1154934000, 1154937600, 1154941200, 1154944800, 
    1154948400, 1154952000, 1154955600, 1154959200, 1154962800, 1154966400, 
    1154970000, 1154973600, 1154977200, 1154980800, 1154984400, 1154988000, 
    1154991600, 1154995200, 1154998800, 1155002400, 1155006000, 1155009600, 
    1155013200, 1155016800, 1155020400, 1155024000, 1155027600, 1155031200, 
    1155034800, 1155038400, 1155042000, 1155045600, 1155049200, 1155052800, 
    1155056400, 1155060000, 1155063600, 1155067200, 1155070800, 1155074400, 
    1155078000, 1155081600, 1155085200, 1155088800, 1155092400, 1155096000, 
    1155099600, 1155103200, 1155106800, 1155110400, 1155114000, 1155117600, 
    1155121200, 1155124800, 1155128400, 1155132000, 1155135600, 1155139200, 
    1155142800, 1155146400, 1155150000, 1155153600, 1155157200, 1155160800, 
    1155164400, 1155168000, 1155171600, 1155175200, 1155178800, 1155182400, 
    1155186000, 1155189600, 1155193200, 1155196800, 1155200400, 1155204000, 
    1155207600, 1155211200, 1155214800, 1155218400, 1155222000, 1155225600, 
    1155229200, 1155232800, 1155236400, 1155240000, 1155243600, 1155247200, 
    1155250800, 1155254400, 1155258000, 1155261600, 1155265200, 1155268800, 
    1155272400, 1155276000, 1155279600, 1155283200, 1155286800, 1155290400, 
    1155294000, 1155297600, 1155301200, 1155304800, 1155308400, 1155312000, 
    1155315600, 1155319200, 1155322800, 1155326400, 1155330000, 1155333600, 
    1155337200, 1155340800, 1155344400, 1155348000, 1155351600, 1155355200, 
    1155358800, 1155362400, 1155366000, 1155369600, 1155373200, 1155376800, 
    1155380400, 1155384000, 1155387600, 1155391200, 1155394800, 1155398400, 
    1155402000, 1155405600, 1155409200, 1155412800, 1155416400, 1155420000, 
    1155423600, 1155427200, 1155430800, 1155434400, 1155438000, 1155441600, 
    1155445200, 1155448800, 1155452400, 1155456000, 1155459600, 1155463200, 
    1155466800, 1155470400, 1155474000, 1155477600, 1155481200, 1155484800, 
    1155488400, 1155492000, 1155495600, 1155499200, 1155502800, 1155506400, 
    1155510000, 1155513600, 1155517200, 1155520800, 1155524400, 1155528000, 
    1155531600, 1155535200, 1155538800, 1155542400, 1155546000, 1155549600, 
    1155553200, 1155556800, 1155560400, 1155564000, 1155567600, 1155571200, 
    1155574800, 1155578400, 1155582000, 1155585600, 1155589200, 1155592800, 
    1155596400, 1155600000, 1155603600, 1155607200, 1155610800, 1155614400, 
    1155618000, 1155621600, 1155625200, 1155628800, 1155632400, 1155636000, 
    1155639600, 1155643200, 1155646800, 1155650400, 1155654000, 1155657600, 
    1155661200, 1155664800, 1155668400, 1155672000, 1155675600, 1155679200, 
    1155682800, 1155686400, 1155690000, 1155693600, 1155697200, 1155700800, 
    1155704400, 1155708000, 1155711600, 1155715200, 1155718800, 1155722400, 
    1155726000, 1155729600, 1155733200, 1155736800, 1155740400, 1155744000, 
    1155747600, 1155751200, 1155754800, 1155758400, 1155762000, 1155765600, 
    1155769200, 1155772800, 1155776400, 1155780000, 1155783600, 1155787200, 
    1155790800, 1155794400, 1155798000, 1155801600, 1155805200, 1155808800, 
    1155812400, 1155816000, 1155819600, 1155823200, 1155826800, 1155830400, 
    1155834000, 1155837600, 1155841200, 1155844800, 1155848400, 1155852000, 
    1155855600, 1155859200, 1155862800, 1155866400, 1155870000, 1155873600, 
    1155877200, 1155880800, 1155884400, 1155888000, 1155891600, 1155895200, 
    1155898800, 1155902400, 1155906000, 1155909600, 1155913200, 1155916800, 
    1155920400, 1155924000, 1155927600, 1155931200, 1155934800, 1155938400, 
    1155942000, 1155945600, 1155949200, 1155952800, 1155956400, 1155960000, 
    1155963600, 1155967200, 1155970800, 1155974400, 1155978000, 1155981600, 
    1155985200, 1155988800, 1155992400, 1155996000, 1155999600, 1156003200, 
    1156006800, 1156010400, 1156014000, 1156017600, 1156021200, 1156024800, 
    1156028400, 1156032000, 1156035600, 1156039200, 1156042800, 1156046400, 
    1156050000, 1156053600, 1156057200, 1156060800, 1156064400, 1156068000, 
    1156071600, 1156075200, 1156078800, 1156082400, 1156086000, 1156089600, 
    1156093200, 1156096800, 1156100400, 1156104000, 1156107600, 1156111200, 
    1156114800, 1156118400, 1156122000, 1156125600, 1156129200, 1156132800, 
    1156136400, 1156140000, 1156143600, 1156147200, 1156150800, 1156154400, 
    1156158000, 1156161600, 1156165200, 1156168800, 1156172400, 1156176000, 
    1156179600, 1156183200, 1156186800, 1156190400, 1156194000, 1156197600, 
    1156201200, 1156204800, 1156208400, 1156212000, 1156215600, 1156219200, 
    1156222800, 1156226400, 1156230000, 1156233600, 1156237200, 1156240800, 
    1156244400, 1156248000, 1156251600, 1156255200, 1156258800, 1156262400, 
    1156266000, 1156269600, 1156273200, 1156276800, 1156280400, 1156284000, 
    1156287600, 1156291200, 1156294800, 1156298400, 1156302000, 1156305600, 
    1156309200, 1156312800, 1156316400, 1156320000, 1156323600, 1156327200, 
    1156330800, 1156334400, 1156338000, 1156341600, 1156345200, 1156348800, 
    1156352400, 1156356000, 1156359600, 1156363200, 1156366800, 1156370400, 
    1156374000, 1156377600, 1156381200, 1156384800, 1156388400, 1156392000, 
    1156395600, 1156399200, 1156402800, 1156406400, 1156410000, 1156413600, 
    1156417200, 1156420800, 1156424400, 1156428000, 1156431600, 1156435200, 
    1156438800, 1156442400, 1156446000, 1156449600, 1156453200, 1156456800, 
    1156460400, 1156464000, 1156467600, 1156471200, 1156474800, 1156478400, 
    1156482000, 1156485600, 1156489200, 1156492800, 1156496400, 1156500000, 
    1156503600, 1156507200, 1156510800, 1156514400, 1156518000, 1156521600, 
    1156525200, 1156528800, 1156532400, 1156536000, 1156539600, 1156543200, 
    1156546800, 1156550400, 1156554000, 1156557600, 1156561200, 1156564800, 
    1156568400, 1156572000, 1156575600, 1156579200, 1156582800, 1156586400, 
    1156590000, 1156593600, 1156597200, 1156600800, 1156604400, 1156608000, 
    1156611600, 1156615200, 1156618800, 1156622400, 1156626000, 1156629600, 
    1156633200, 1156636800, 1156640400, 1156644000, 1156647600, 1156651200, 
    1156654800, 1156658400, 1156662000, 1156665600, 1156669200, 1156672800, 
    1156676400, 1156680000, 1156683600, 1156687200, 1156690800, 1156694400, 
    1156698000, 1156701600, 1156705200, 1156708800, 1156712400, 1156716000, 
    1156719600, 1156723200, 1156726800, 1156730400, 1156734000, 1156737600, 
    1156741200, 1156744800, 1156748400, 1156752000, 1156755600, 1156759200, 
    1156762800, 1156766400, 1156770000, 1156773600, 1156777200, 1156780800, 
    1156784400, 1156788000, 1156791600, 1156795200, 1156798800, 1156802400, 
    1156806000, 1156809600, 1156813200, 1156816800, 1156820400, 1156824000, 
    1156827600, 1156831200, 1156834800, 1156838400, 1156842000, 1156845600, 
    1156849200, 1156852800, 1156856400, 1156860000, 1156863600, 1156867200, 
    1156870800, 1156874400, 1156878000, 1156881600, 1156885200, 1156888800, 
    1156892400, 1156896000, 1156899600, 1156903200, 1156906800, 1156910400, 
    1156914000, 1156917600, 1156921200, 1156924800, 1156928400, 1156932000, 
    1156935600, 1156939200, 1156942800, 1156946400, 1156950000, 1156953600, 
    1156957200, 1156960800, 1156964400, 1156968000, 1156971600, 1156975200, 
    1156978800, 1156982400, 1156986000, 1156989600, 1156993200, 1156996800, 
    1157000400, 1157004000, 1157007600, 1157011200, 1157014800, 1157018400, 
    1157022000, 1157025600, 1157029200, 1157032800, 1157036400, 1157040000, 
    1157043600, 1157047200, 1157050800, 1157054400, 1157058000, 1157061600, 
    1157065200, 1157068800, 1157072400, 1157076000, 1157079600, 1157083200, 
    1157086800, 1157090400, 1157094000, 1157097600, 1157101200, 1157104800, 
    1157108400, 1157112000, 1157115600, 1157119200, 1157122800, 1157126400, 
    1157130000, 1157133600, 1157137200, 1157140800, 1157144400, 1157148000, 
    1157151600, 1157155200, 1157158800, 1157162400, 1157166000, 1157169600, 
    1157173200, 1157176800, 1157180400, 1157184000, 1157187600, 1157191200, 
    1157194800, 1157198400, 1157202000, 1157205600, 1157209200, 1157212800, 
    1157216400, 1157220000, 1157223600, 1157227200, 1157230800, 1157234400, 
    1157238000, 1157241600, 1157245200, 1157248800, 1157252400, 1157256000, 
    1157259600, 1157263200, 1157266800, 1157270400, 1157274000, 1157277600, 
    1157281200, 1157284800, 1157288400, 1157292000, 1157295600, 1157299200, 
    1157302800, 1157306400, 1157310000, 1157313600, 1157317200, 1157320800, 
    1157324400, 1157328000, 1157331600, 1157335200, 1157338800, 1157342400, 
    1157346000, 1157349600, 1157353200, 1157356800, 1157360400, 1157364000, 
    1157367600, 1157371200, 1157374800, 1157378400, 1157382000, 1157385600, 
    1157389200, 1157392800, 1157396400, 1157400000, 1157403600, 1157407200, 
    1157410800, 1157414400, 1157418000, 1157421600, 1157425200, 1157428800, 
    1157432400, 1157436000, 1157439600, 1157443200, 1157446800, 1157450400, 
    1157454000, 1157457600, 1157461200, 1157464800, 1157468400, 1157472000, 
    1157475600, 1157479200, 1157482800, 1157486400, 1157490000, 1157493600, 
    1157497200, 1157500800, 1157504400, 1157508000, 1157511600, 1157515200, 
    1157518800, 1157522400, 1157526000, 1157529600, 1157533200, 1157536800, 
    1157540400, 1157544000, 1157547600, 1157551200, 1157554800, 1157558400, 
    1157562000, 1157565600, 1157569200, 1157572800, 1157576400, 1157580000, 
    1157583600, 1157587200, 1157590800, 1157594400, 1157598000, 1157601600, 
    1157605200, 1157608800, 1157612400, 1157616000, 1157619600, 1157623200, 
    1157626800, 1157630400, 1157634000, 1157637600, 1157641200, 1157644800, 
    1157648400, 1157652000, 1157655600, 1157659200, 1157662800, 1157666400, 
    1157670000, 1157673600, 1157677200, 1157680800, 1157684400, 1157688000, 
    1157691600, 1157695200, 1157698800, 1157702400, 1157706000, 1157709600, 
    1157713200, 1157716800, 1157720400, 1157724000, 1157727600, 1157731200, 
    1157734800, 1157738400, 1157742000, 1157745600, 1157749200, 1157752800, 
    1157756400, 1157760000, 1157763600, 1157767200, 1157770800, 1157774400, 
    1157778000, 1157781600, 1157785200, 1157788800, 1157792400, 1157796000, 
    1157799600, 1157803200, 1157806800, 1157810400, 1157814000, 1157817600, 
    1157821200, 1157824800, 1157828400, 1157832000, 1157835600, 1157839200, 
    1157842800, 1157846400, 1157850000, 1157853600, 1157857200, 1157860800, 
    1157864400, 1157868000, 1157871600, 1157875200, 1157878800, 1157882400, 
    1157886000, 1157889600, 1157893200, 1157896800, 1157900400, 1157904000, 
    1157907600, 1157911200, 1157914800, 1157918400, 1157922000, 1157925600, 
    1157929200, 1157932800, 1157936400, 1157940000, 1157943600, 1157947200, 
    1157950800, 1157954400, 1157958000, 1157961600, 1157965200, 1157968800, 
    1157972400, 1157976000, 1157979600, 1157983200, 1157986800, 1157990400, 
    1157994000, 1157997600, 1158001200, 1158004800, 1158008400, 1158012000, 
    1158015600, 1158019200, 1158022800, 1158026400, 1158030000, 1158033600, 
    1158037200, 1158040800, 1158044400, 1158048000, 1158051600, 1158055200, 
    1158058800, 1158062400, 1158066000, 1158069600, 1158073200, 1158076800, 
    1158080400, 1158084000, 1158087600, 1158091200, 1158094800, 1158098400, 
    1158102000, 1158105600, 1158109200, 1158112800, 1158116400, 1158120000, 
    1158123600, 1158127200, 1158130800, 1158134400, 1158138000, 1158141600, 
    1158145200, 1158148800, 1158152400, 1158156000, 1158159600, 1158163200, 
    1158166800, 1158170400, 1158174000, 1158177600, 1158181200, 1158184800, 
    1158188400, 1158192000, 1158195600, 1158199200, 1158202800, 1158206400, 
    1158210000, 1158213600, 1158217200, 1158220800, 1158224400, 1158228000, 
    1158231600, 1158235200, 1158238800, 1158242400, 1158246000, 1158249600, 
    1158253200, 1158256800, 1158260400, 1158264000, 1158267600, 1158271200, 
    1158274800, 1158278400, 1158282000, 1158285600, 1158289200, 1158292800, 
    1158296400, 1158300000, 1158303600, 1158307200, 1158310800, 1158314400, 
    1158318000, 1158321600, 1158325200, 1158328800, 1158332400, 1158336000, 
    1158339600, 1158343200, 1158346800, 1158350400, 1158354000, 1158357600, 
    1158361200, 1158364800, 1158368400, 1158372000, 1158375600, 1158379200, 
    1158382800, 1158386400, 1158390000, 1158393600, 1158397200, 1158400800, 
    1158404400, 1158408000, 1158411600, 1158415200, 1158418800, 1158422400, 
    1158426000, 1158429600, 1158433200, 1158436800, 1158440400, 1158444000, 
    1158447600, 1158451200, 1158454800, 1158458400, 1158462000, 1158465600, 
    1158469200, 1158472800, 1158476400, 1158480000, 1158483600, 1158487200, 
    1158490800, 1158494400, 1158498000, 1158501600, 1158505200, 1158508800, 
    1158512400, 1158516000, 1158519600, 1158523200, 1158526800, 1158530400, 
    1158534000, 1158537600, 1158541200, 1158544800, 1158548400, 1158552000, 
    1158555600, 1158559200, 1158562800, 1158566400, 1158570000, 1158573600, 
    1158577200, 1158580800, 1158584400, 1158588000, 1158591600, 1158595200, 
    1158598800, 1158602400, 1158606000, 1158609600, 1158613200, 1158616800, 
    1158620400, 1158624000, 1158627600, 1158631200, 1158634800, 1158638400, 
    1158642000, 1158645600, 1158649200, 1158652800, 1158656400, 1158660000, 
    1158663600, 1158667200, 1158670800, 1158674400, 1158678000, 1158681600, 
    1158685200, 1158688800, 1158692400, 1158696000, 1158699600, 1158703200, 
    1158706800, 1158710400, 1158714000, 1158717600, 1158721200, 1158724800, 
    1158728400, 1158732000, 1158735600, 1158739200, 1158742800, 1158746400, 
    1158750000, 1158753600, 1158757200, 1158760800, 1158764400, 1158768000, 
    1158771600, 1158775200, 1158778800, 1158782400, 1158786000, 1158789600, 
    1158793200, 1158796800, 1158800400, 1158804000, 1158807600, 1158811200, 
    1158814800, 1158818400, 1158822000, 1158825600, 1158829200, 1158832800, 
    1158836400, 1158840000, 1158843600, 1158847200, 1158850800, 1158854400, 
    1158858000, 1158861600, 1158865200, 1158868800, 1158872400, 1158876000, 
    1158879600, 1158883200, 1158886800, 1158890400, 1158894000, 1158897600, 
    1158901200, 1158904800, 1158908400, 1158912000, 1158915600, 1158919200, 
    1158922800, 1158926400, 1158930000, 1158933600, 1158937200, 1158940800, 
    1158944400, 1158948000, 1158951600, 1158955200, 1158958800, 1158962400, 
    1158966000, 1158969600, 1158973200, 1158976800, 1158980400, 1158984000, 
    1158987600, 1158991200, 1158994800, 1158998400, 1159002000, 1159005600, 
    1159009200, 1159012800, 1159016400, 1159020000, 1159023600, 1159027200, 
    1159030800, 1159034400, 1159038000, 1159041600, 1159045200, 1159048800, 
    1159052400, 1159056000, 1159059600, 1159063200, 1159066800, 1159070400, 
    1159074000, 1159077600, 1159081200, 1159084800, 1159088400, 1159092000, 
    1159095600, 1159099200, 1159102800, 1159106400, 1159110000, 1159113600, 
    1159117200, 1159120800, 1159124400, 1159128000, 1159131600, 1159135200, 
    1159138800, 1159142400, 1159146000, 1159149600, 1159153200, 1159156800, 
    1159160400, 1159164000, 1159167600, 1159171200, 1159174800, 1159178400, 
    1159182000, 1159185600, 1159189200, 1159192800, 1159196400, 1159200000, 
    1159203600, 1159207200, 1159210800, 1159214400, 1159218000, 1159221600, 
    1159225200, 1159228800, 1159232400, 1159236000, 1159239600, 1159243200, 
    1159246800, 1159250400, 1159254000, 1159257600, 1159261200, 1159264800, 
    1159268400, 1159272000, 1159275600, 1159279200, 1159282800, 1159286400, 
    1159290000, 1159293600, 1159297200, 1159300800, 1159304400, 1159308000, 
    1159311600, 1159315200, 1159318800, 1159322400, 1159326000, 1159329600, 
    1159333200, 1159336800, 1159340400, 1159344000, 1159347600, 1159351200, 
    1159354800, 1159358400, 1159362000, 1159365600, 1159369200, 1159372800, 
    1159376400, 1159380000, 1159383600, 1159387200, 1159390800, 1159394400, 
    1159398000, 1159401600, 1159405200, 1159408800, 1159412400, 1159416000, 
    1159419600, 1159423200, 1159426800, 1159430400, 1159434000, 1159437600, 
    1159441200, 1159444800, 1159448400, 1159452000, 1159455600, 1159459200, 
    1159462800, 1159466400, 1159470000, 1159473600, 1159477200, 1159480800, 
    1159484400, 1159488000, 1159491600, 1159495200, 1159498800, 1159502400, 
    1159506000, 1159509600, 1159513200, 1159516800, 1159520400, 1159524000, 
    1159527600, 1159531200, 1159534800, 1159538400, 1159542000, 1159545600, 
    1159549200, 1159552800, 1159556400, 1159560000, 1159563600, 1159567200, 
    1159570800, 1159574400, 1159578000, 1159581600, 1159585200, 1159588800, 
    1159592400, 1159596000, 1159599600, 1159603200, 1159606800, 1159610400, 
    1159614000, 1159617600, 1159621200, 1159624800, 1159628400, 1159632000, 
    1159635600, 1159639200, 1159642800, 1159646400, 1159650000, 1159653600, 
    1159657200, 1159660800, 1159664400, 1159668000, 1159671600, 1159675200, 
    1159678800, 1159682400, 1159686000, 1159689600, 1159693200, 1159696800, 
    1159700400, 1159704000, 1159707600, 1159711200, 1159714800, 1159718400, 
    1159722000, 1159725600, 1159729200, 1159732800, 1159736400, 1159740000, 
    1159743600, 1159747200, 1159750800, 1159754400, 1159758000, 1159761600, 
    1159765200, 1159768800, 1159772400, 1159776000, 1159779600, 1159783200, 
    1159786800, 1159790400, 1159794000, 1159797600, 1159801200, 1159804800, 
    1159808400, 1159812000, 1159815600, 1159819200, 1159822800, 1159826400, 
    1159830000, 1159833600, 1159837200, 1159840800, 1159844400, 1159848000, 
    1159851600, 1159855200, 1159858800, 1159862400, 1159866000, 1159869600, 
    1159873200, 1159876800, 1159880400, 1159884000, 1159887600, 1159891200, 
    1159894800, 1159898400, 1159902000, 1159905600, 1159909200, 1159912800, 
    1159916400, 1159920000, 1159923600, 1159927200, 1159930800, 1159934400, 
    1159938000, 1159941600, 1159945200, 1159948800, 1159952400, 1159956000, 
    1159959600, 1159963200, 1159966800, 1159970400, 1159974000, 1159977600, 
    1159981200, 1159984800, 1159988400, 1159992000, 1159995600, 1159999200, 
    1160002800, 1160006400, 1160010000, 1160013600, 1160017200, 1160020800, 
    1160024400, 1160028000, 1160031600, 1160035200, 1160038800, 1160042400, 
    1160046000, 1160049600, 1160053200, 1160056800, 1160060400, 1160064000, 
    1160067600, 1160071200, 1160074800, 1160078400, 1160082000, 1160085600, 
    1160089200, 1160092800, 1160096400, 1160100000, 1160103600, 1160107200, 
    1160110800, 1160114400, 1160118000, 1160121600, 1160125200, 1160128800, 
    1160132400, 1160136000, 1160139600, 1160143200, 1160146800, 1160150400, 
    1160154000, 1160157600, 1160161200, 1160164800, 1160168400, 1160172000, 
    1160175600, 1160179200, 1160182800, 1160186400, 1160190000, 1160193600, 
    1160197200, 1160200800, 1160204400, 1160208000, 1160211600, 1160215200, 
    1160218800, 1160222400, 1160226000, 1160229600, 1160233200, 1160236800, 
    1160240400, 1160244000, 1160247600, 1160251200, 1160254800, 1160258400, 
    1160262000, 1160265600, 1160269200, 1160272800, 1160276400, 1160280000, 
    1160283600, 1160287200, 1160290800, 1160294400, 1160298000, 1160301600, 
    1160305200, 1160308800, 1160312400, 1160316000, 1160319600, 1160323200, 
    1160326800, 1160330400, 1160334000, 1160337600, 1160341200, 1160344800, 
    1160348400, 1160352000, 1160355600, 1160359200, 1160362800, 1160366400, 
    1160370000, 1160373600, 1160377200, 1160380800, 1160384400, 1160388000, 
    1160391600, 1160395200, 1160398800, 1160402400, 1160406000, 1160409600, 
    1160413200, 1160416800, 1160420400, 1160424000, 1160427600, 1160431200, 
    1160434800, 1160438400, 1160442000, 1160445600, 1160449200, 1160452800, 
    1160456400, 1160460000, 1160463600, 1160467200, 1160470800, 1160474400, 
    1160478000, 1160481600, 1160485200, 1160488800, 1160492400, 1160496000, 
    1160499600, 1160503200, 1160506800, 1160510400, 1160514000, 1160517600, 
    1160521200, 1160524800, 1160528400, 1160532000, 1160535600, 1160539200, 
    1160542800, 1160546400, 1160550000, 1160553600, 1160557200, 1160560800, 
    1160564400, 1160568000, 1160571600, 1160575200, 1160578800, 1160582400, 
    1160586000, 1160589600, 1160593200, 1160596800, 1160600400, 1160604000, 
    1160607600, 1160611200, 1160614800, 1160618400, 1160622000, 1160625600, 
    1160629200, 1160632800, 1160636400, 1160640000, 1160643600, 1160647200, 
    1160650800, 1160654400, 1160658000, 1160661600, 1160665200, 1160668800, 
    1160672400, 1160676000, 1160679600, 1160683200, 1160686800, 1160690400, 
    1160694000, 1160697600, 1160701200, 1160704800, 1160708400, 1160712000, 
    1160715600, 1160719200, 1160722800, 1160726400, 1160730000, 1160733600, 
    1160737200, 1160740800, 1160744400, 1160748000, 1160751600, 1160755200, 
    1160758800, 1160762400, 1160766000, 1160769600, 1160773200, 1160776800, 
    1160780400, 1160784000, 1160787600, 1160791200, 1160794800, 1160798400, 
    1160802000, 1160805600, 1160809200, 1160812800, 1160816400, 1160820000, 
    1160823600, 1160827200, 1160830800, 1160834400, 1160838000, 1160841600, 
    1160845200, 1160848800, 1160852400, 1160856000, 1160859600, 1160863200, 
    1160866800, 1160870400, 1160874000, 1160877600, 1160881200, 1160884800, 
    1160888400, 1160892000, 1160895600, 1160899200, 1160902800, 1160906400, 
    1160910000, 1160913600, 1160917200, 1160920800, 1160924400, 1160928000, 
    1160931600, 1160935200, 1160938800, 1160942400, 1160946000, 1160949600, 
    1160953200, 1160956800, 1160960400, 1160964000, 1160967600, 1160971200, 
    1160974800, 1160978400, 1160982000, 1160985600, 1160989200, 1160992800, 
    1160996400, 1161000000, 1161003600, 1161007200, 1161010800, 1161014400, 
    1161018000, 1161021600, 1161025200, 1161028800, 1161032400, 1161036000, 
    1161039600, 1161043200, 1161046800, 1161050400, 1161054000, 1161057600, 
    1161061200, 1161064800, 1161068400, 1161072000, 1161075600, 1161079200, 
    1161082800, 1161086400, 1161090000, 1161093600, 1161097200, 1161100800, 
    1161104400, 1161108000, 1161111600, 1161115200, 1161118800, 1161122400, 
    1161126000, 1161129600, 1161133200, 1161136800, 1161140400, 1161144000, 
    1161147600, 1161151200, 1161154800, 1161158400, 1161162000, 1161165600, 
    1161169200, 1161172800, 1161176400, 1161180000, 1161183600, 1161187200, 
    1161190800, 1161194400, 1161198000, 1161201600, 1161205200, 1161208800, 
    1161212400, 1161216000, 1161219600, 1161223200, 1161226800, 1161230400, 
    1161234000, 1161237600, 1161241200, 1161244800, 1161248400, 1161252000, 
    1161255600, 1161259200, 1161262800, 1161266400, 1161270000, 1161273600, 
    1161277200, 1161280800, 1161284400, 1161288000, 1161291600, 1161295200, 
    1161298800, 1161302400, 1161306000, 1161309600, 1161313200, 1161316800, 
    1161320400, 1161324000, 1161327600, 1161331200, 1161334800, 1161338400, 
    1161342000, 1161345600, 1161349200, 1161352800, 1161356400, 1161360000, 
    1161363600, 1161367200, 1161370800, 1161374400, 1161378000, 1161381600, 
    1161385200, 1161388800, 1161392400, 1161396000, 1161399600, 1161403200, 
    1161406800, 1161410400, 1161414000, 1161417600, 1161421200, 1161424800, 
    1161428400, 1161432000, 1161435600, 1161439200, 1161442800, 1161446400, 
    1161450000, 1161453600, 1161457200, 1161460800, 1161464400, 1161468000, 
    1161471600, 1161475200, 1161478800, 1161482400, 1161486000, 1161489600, 
    1161493200, 1161496800, 1161500400, 1161504000, 1161507600, 1161511200, 
    1161514800, 1161518400, 1161522000, 1161525600, 1161529200, 1161532800, 
    1161536400, 1161540000, 1161543600, 1161547200, 1161550800, 1161554400, 
    1161558000, 1161561600, 1161565200, 1161568800, 1161572400, 1161576000, 
    1161579600, 1161583200, 1161586800, 1161590400, 1161594000, 1161597600, 
    1161601200, 1161604800, 1161608400, 1161612000, 1161615600, 1161619200, 
    1161622800, 1161626400, 1161630000, 1161633600, 1161637200, 1161640800, 
    1161644400, 1161648000, 1161651600, 1161655200, 1161658800, 1161662400, 
    1161666000, 1161669600, 1161673200, 1161676800, 1161680400, 1161684000, 
    1161687600, 1161691200, 1161694800, 1161698400, 1161702000, 1161705600, 
    1161709200, 1161712800, 1161716400, 1161720000, 1161723600, 1161727200, 
    1161730800, 1161734400, 1161738000, 1161741600, 1161745200, 1161748800, 
    1161752400, 1161756000, 1161759600, 1161763200, 1161766800, 1161770400, 
    1161774000, 1161777600, 1161781200, 1161784800, 1161788400, 1161792000, 
    1161795600, 1161799200, 1161802800, 1161806400, 1161810000, 1161813600, 
    1161817200, 1161820800, 1161824400, 1161828000, 1161831600, 1161835200, 
    1161838800, 1161842400, 1161846000, 1161849600, 1161853200, 1161856800, 
    1161860400, 1161864000, 1161867600, 1161871200, 1161874800, 1161878400, 
    1161882000, 1161885600, 1161889200, 1161892800, 1161896400, 1161900000, 
    1161903600, 1161907200, 1161910800, 1161914400, 1161918000, 1161921600, 
    1161925200, 1161928800, 1161932400, 1161936000, 1161939600, 1161943200, 
    1161946800, 1161950400, 1161954000, 1161957600, 1161961200, 1161964800, 
    1161968400, 1161972000, 1161975600, 1161979200, 1161982800, 1161986400, 
    1161990000, 1161993600, 1161997200, 1162000800, 1162004400, 1162008000, 
    1162011600, 1162015200, 1162018800, 1162022400, 1162026000, 1162029600, 
    1162033200, 1162036800, 1162040400, 1162044000, 1162047600, 1162051200, 
    1162054800, 1162058400, 1162062000, 1162065600, 1162069200, 1162072800, 
    1162076400, 1162080000, 1162083600, 1162087200, 1162090800, 1162094400, 
    1162098000, 1162101600, 1162105200, 1162108800, 1162112400, 1162116000, 
    1162119600, 1162123200, 1162126800, 1162130400, 1162134000, 1162137600, 
    1162141200, 1162144800, 1162148400, 1162152000, 1162155600, 1162159200, 
    1162162800, 1162166400, 1162170000, 1162173600, 1162177200, 1162180800, 
    1162184400, 1162188000, 1162191600, 1162195200, 1162198800, 1162202400, 
    1162206000, 1162209600, 1162213200, 1162216800, 1162220400, 1162224000, 
    1162227600, 1162231200, 1162234800, 1162238400, 1162242000, 1162245600, 
    1162249200, 1162252800, 1162256400, 1162260000, 1162263600, 1162267200, 
    1162270800, 1162274400, 1162278000, 1162281600, 1162285200, 1162288800, 
    1162292400, 1162296000, 1162299600, 1162303200, 1162306800, 1162310400, 
    1162314000, 1162317600, 1162321200, 1162324800, 1162328400, 1162332000, 
    1162335600, 1162339200, 1162342800, 1162346400, 1162350000, 1162353600, 
    1162357200, 1162360800, 1162364400, 1162368000, 1162371600, 1162375200, 
    1162378800, 1162382400, 1162386000, 1162389600, 1162393200, 1162396800, 
    1162400400, 1162404000, 1162407600, 1162411200, 1162414800, 1162418400, 
    1162422000, 1162425600, 1162429200, 1162432800, 1162436400, 1162440000, 
    1162443600, 1162447200, 1162450800, 1162454400, 1162458000, 1162461600, 
    1162465200, 1162468800, 1162472400, 1162476000, 1162479600, 1162483200, 
    1162486800, 1162490400, 1162494000, 1162497600, 1162501200, 1162504800, 
    1162508400, 1162512000, 1162515600, 1162519200, 1162522800, 1162526400, 
    1162530000, 1162533600, 1162537200, 1162540800, 1162544400, 1162548000, 
    1162551600, 1162555200, 1162558800, 1162562400, 1162566000, 1162569600, 
    1162573200, 1162576800, 1162580400, 1162584000, 1162587600, 1162591200, 
    1162594800, 1162598400, 1162602000, 1162605600, 1162609200, 1162612800, 
    1162616400, 1162620000, 1162623600, 1162627200, 1162630800, 1162634400, 
    1162638000, 1162641600, 1162645200, 1162648800, 1162652400, 1162656000, 
    1162659600, 1162663200, 1162666800, 1162670400, 1162674000, 1162677600, 
    1162681200, 1162684800, 1162688400, 1162692000, 1162695600, 1162699200, 
    1162702800, 1162706400, 1162710000, 1162713600, 1162717200, 1162720800, 
    1162724400, 1162728000, 1162731600, 1162735200, 1162738800, 1162742400, 
    1162746000, 1162749600, 1162753200, 1162756800, 1162760400, 1162764000, 
    1162767600, 1162771200, 1162774800, 1162778400, 1162782000, 1162785600, 
    1162789200, 1162792800, 1162796400, 1162800000, 1162803600, 1162807200, 
    1162810800, 1162814400, 1162818000, 1162821600, 1162825200, 1162828800, 
    1162832400, 1162836000, 1162839600, 1162843200, 1162846800, 1162850400, 
    1162854000, 1162857600, 1162861200, 1162864800, 1162868400, 1162872000, 
    1162875600, 1162879200, 1162882800, 1162886400, 1162890000, 1162893600, 
    1162897200, 1162900800, 1162904400, 1162908000, 1162911600, 1162915200, 
    1162918800, 1162922400, 1162926000, 1162929600, 1162933200, 1162936800, 
    1162940400, 1162944000, 1162947600, 1162951200, 1162954800, 1162958400, 
    1162962000, 1162965600, 1162969200, 1162972800, 1162976400, 1162980000, 
    1162983600, 1162987200, 1162990800, 1162994400, 1162998000, 1163001600, 
    1163005200, 1163008800, 1163012400, 1163016000, 1163019600, 1163023200, 
    1163026800, 1163030400, 1163034000, 1163037600, 1163041200, 1163044800, 
    1163048400, 1163052000, 1163055600, 1163059200, 1163062800, 1163066400, 
    1163070000, 1163073600, 1163077200, 1163080800, 1163084400, 1163088000, 
    1163091600, 1163095200, 1163098800, 1163102400, 1163106000, 1163109600, 
    1163113200, 1163116800, 1163120400, 1163124000, 1163127600, 1163131200, 
    1163134800, 1163138400, 1163142000, 1163145600, 1163149200, 1163152800, 
    1163156400, 1163160000, 1163163600, 1163167200, 1163170800, 1163174400, 
    1163178000, 1163181600, 1163185200, 1163188800, 1163192400, 1163196000, 
    1163199600, 1163203200, 1163206800, 1163210400, 1163214000, 1163217600, 
    1163221200, 1163224800, 1163228400, 1163232000, 1163235600, 1163239200, 
    1163242800, 1163246400, 1163250000, 1163253600, 1163257200, 1163260800, 
    1163264400, 1163268000, 1163271600, 1163275200, 1163278800, 1163282400, 
    1163286000, 1163289600, 1163293200, 1163296800, 1163300400, 1163304000, 
    1163307600, 1163311200, 1163314800, 1163318400, 1163322000, 1163325600, 
    1163329200, 1163332800, 1163336400, 1163340000, 1163343600, 1163347200, 
    1163350800, 1163354400, 1163358000, 1163361600, 1163365200, 1163368800, 
    1163372400, 1163376000, 1163379600, 1163383200, 1163386800, 1163390400, 
    1163394000, 1163397600, 1163401200, 1163404800, 1163408400, 1163412000, 
    1163415600, 1163419200, 1163422800, 1163426400, 1163430000, 1163433600, 
    1163437200, 1163440800, 1163444400, 1163448000, 1163451600, 1163455200, 
    1163458800, 1163462400, 1163466000, 1163469600, 1163473200, 1163476800, 
    1163480400, 1163484000, 1163487600, 1163491200, 1163494800, 1163498400, 
    1163502000, 1163505600, 1163509200, 1163512800, 1163516400, 1163520000, 
    1163523600, 1163527200, 1163530800, 1163534400, 1163538000, 1163541600, 
    1163545200, 1163548800, 1163552400, 1163556000, 1163559600, 1163563200, 
    1163566800, 1163570400, 1163574000, 1163577600, 1163581200, 1163584800, 
    1163588400, 1163592000, 1163595600, 1163599200, 1163602800, 1163606400, 
    1163610000, 1163613600, 1163617200, 1163620800, 1163624400, 1163628000, 
    1163631600, 1163635200, 1163638800, 1163642400, 1163646000, 1163649600, 
    1163653200, 1163656800, 1163660400, 1163664000, 1163667600, 1163671200, 
    1163674800, 1163678400, 1163682000, 1163685600, 1163689200, 1163692800, 
    1163696400, 1163700000, 1163703600, 1163707200, 1163710800, 1163714400, 
    1163718000, 1163721600, 1163725200, 1163728800, 1163732400, 1163736000, 
    1163739600, 1163743200, 1163746800, 1163750400, 1163754000, 1163757600, 
    1163761200, 1163764800, 1163768400, 1163772000, 1163775600, 1163779200, 
    1163782800, 1163786400, 1163790000, 1163793600, 1163797200, 1163800800, 
    1163804400, 1163808000, 1163811600, 1163815200, 1163818800, 1163822400, 
    1163826000, 1163829600, 1163833200, 1163836800, 1163840400, 1163844000, 
    1163847600, 1163851200, 1163854800, 1163858400, 1163862000, 1163865600, 
    1163869200, 1163872800, 1163876400, 1163880000, 1163883600, 1163887200, 
    1163890800, 1163894400, 1163898000, 1163901600, 1163905200, 1163908800, 
    1163912400, 1163916000, 1163919600, 1163923200, 1163926800, 1163930400, 
    1163934000, 1163937600, 1163941200, 1163944800, 1163948400, 1163952000, 
    1163955600, 1163959200, 1163962800, 1163966400, 1163970000, 1163973600, 
    1163977200, 1163980800, 1163984400, 1163988000, 1163991600, 1163995200, 
    1163998800, 1164002400, 1164006000, 1164009600, 1164013200, 1164016800, 
    1164020400, 1164024000, 1164027600, 1164031200, 1164034800, 1164038400, 
    1164042000, 1164045600, 1164049200, 1164052800, 1164056400, 1164060000, 
    1164063600, 1164067200, 1164070800, 1164074400, 1164078000, 1164081600, 
    1164085200, 1164088800, 1164092400, 1164096000, 1164099600, 1164103200, 
    1164106800, 1164110400, 1164114000, 1164117600, 1164121200, 1164124800, 
    1164128400, 1164132000, 1164135600, 1164139200, 1164142800, 1164146400, 
    1164150000, 1164153600, 1164157200, 1164160800, 1164164400, 1164168000, 
    1164171600, 1164175200, 1164178800, 1164182400, 1164186000, 1164189600, 
    1164193200, 1164196800, 1164200400, 1164204000, 1164207600, 1164211200, 
    1164214800, 1164218400, 1164222000, 1164225600, 1164229200, 1164232800, 
    1164236400, 1164240000, 1164243600, 1164247200, 1164250800, 1164254400, 
    1164258000, 1164261600, 1164265200, 1164268800, 1164272400, 1164276000, 
    1164279600, 1164283200, 1164286800, 1164290400, 1164294000, 1164297600, 
    1164301200, 1164304800, 1164308400, 1164312000, 1164315600, 1164319200, 
    1164322800, 1164326400, 1164330000, 1164333600, 1164337200, 1164340800, 
    1164344400, 1164348000, 1164351600, 1164355200, 1164358800, 1164362400, 
    1164366000, 1164369600, 1164373200, 1164376800, 1164380400, 1164384000, 
    1164387600, 1164391200, 1164394800, 1164398400, 1164402000, 1164405600, 
    1164409200, 1164412800, 1164416400, 1164420000, 1164423600, 1164427200, 
    1164430800, 1164434400, 1164438000, 1164441600, 1164445200, 1164448800, 
    1164452400, 1164456000, 1164459600, 1164463200, 1164466800, 1164470400, 
    1164474000, 1164477600, 1164481200, 1164484800, 1164488400, 1164492000, 
    1164495600, 1164499200, 1164502800, 1164506400, 1164510000, 1164513600, 
    1164517200, 1164520800, 1164524400, 1164528000, 1164531600, 1164535200, 
    1164538800, 1164542400, 1164546000, 1164549600, 1164553200, 1164556800, 
    1164560400, 1164564000, 1164567600, 1164571200, 1164574800, 1164578400, 
    1164582000, 1164585600, 1164589200, 1164592800, 1164596400, 1164600000, 
    1164603600, 1164607200, 1164610800, 1164614400, 1164618000, 1164621600, 
    1164625200, 1164628800, 1164632400, 1164636000, 1164639600, 1164643200, 
    1164646800, 1164650400, 1164654000, 1164657600, 1164661200, 1164664800, 
    1164668400, 1164672000, 1164675600, 1164679200, 1164682800, 1164686400, 
    1164690000, 1164693600, 1164697200, 1164700800, 1164704400, 1164708000, 
    1164711600, 1164715200, 1164718800, 1164722400, 1164726000, 1164729600, 
    1164733200, 1164736800, 1164740400, 1164744000, 1164747600, 1164751200, 
    1164754800, 1164758400, 1164762000, 1164765600, 1164769200, 1164772800, 
    1164776400, 1164780000, 1164783600, 1164787200, 1164790800, 1164794400, 
    1164798000, 1164801600, 1164805200, 1164808800, 1164812400, 1164816000, 
    1164819600, 1164823200, 1164826800, 1164830400, 1164834000, 1164837600, 
    1164841200, 1164844800, 1164848400, 1164852000, 1164855600, 1164859200, 
    1164862800, 1164866400, 1164870000, 1164873600, 1164877200, 1164880800, 
    1164884400, 1164888000, 1164891600, 1164895200, 1164898800, 1164902400, 
    1164906000, 1164909600, 1164913200, 1164916800, 1164920400, 1164924000, 
    1164927600, 1164931200, 1164934800, 1164938400, 1164942000, 1164945600, 
    1164949200, 1164952800, 1164956400, 1164960000, 1164963600, 1164967200, 
    1164970800, 1164974400, 1164978000, 1164981600, 1164985200, 1164988800, 
    1164992400, 1164996000, 1164999600, 1165003200, 1165006800, 1165010400, 
    1165014000, 1165017600, 1165021200, 1165024800, 1165028400, 1165032000, 
    1165035600, 1165039200, 1165042800, 1165046400, 1165050000, 1165053600, 
    1165057200, 1165060800, 1165064400, 1165068000, 1165071600, 1165075200, 
    1165078800, 1165082400, 1165086000, 1165089600, 1165093200, 1165096800, 
    1165100400, 1165104000, 1165107600, 1165111200, 1165114800, 1165118400, 
    1165122000, 1165125600, 1165129200, 1165132800, 1165136400, 1165140000, 
    1165143600, 1165147200, 1165150800, 1165154400, 1165158000, 1165161600, 
    1165165200, 1165168800, 1165172400, 1165176000, 1165179600, 1165183200, 
    1165186800, 1165190400, 1165194000, 1165197600, 1165201200, 1165204800, 
    1165208400, 1165212000, 1165215600, 1165219200, 1165222800, 1165226400, 
    1165230000, 1165233600, 1165237200, 1165240800, 1165244400, 1165248000, 
    1165251600, 1165255200, 1165258800, 1165262400, 1165266000, 1165269600, 
    1165273200, 1165276800, 1165280400, 1165284000, 1165287600, 1165291200, 
    1165294800, 1165298400, 1165302000, 1165305600, 1165309200, 1165312800, 
    1165316400, 1165320000, 1165323600, 1165327200, 1165330800, 1165334400, 
    1165338000, 1165341600, 1165345200, 1165348800, 1165352400, 1165356000, 
    1165359600, 1165363200, 1165366800, 1165370400, 1165374000, 1165377600, 
    1165381200, 1165384800, 1165388400, 1165392000, 1165395600, 1165399200, 
    1165402800, 1165406400, 1165410000, 1165413600, 1165417200, 1165420800, 
    1165424400, 1165428000, 1165431600, 1165435200, 1165438800, 1165442400, 
    1165446000, 1165449600, 1165453200, 1165456800, 1165460400, 1165464000, 
    1165467600, 1165471200, 1165474800, 1165478400, 1165482000, 1165485600, 
    1165489200, 1165492800, 1165496400, 1165500000, 1165503600, 1165507200, 
    1165510800, 1165514400, 1165518000, 1165521600, 1165525200, 1165528800, 
    1165532400, 1165536000, 1165539600, 1165543200, 1165546800, 1165550400, 
    1165554000, 1165557600, 1165561200, 1165564800, 1165568400, 1165572000, 
    1165575600, 1165579200, 1165582800, 1165586400, 1165590000, 1165593600, 
    1165597200, 1165600800, 1165604400, 1165608000, 1165611600, 1165615200, 
    1165618800, 1165622400, 1165626000, 1165629600, 1165633200, 1165636800, 
    1165640400, 1165644000, 1165647600, 1165651200, 1165654800, 1165658400, 
    1165662000, 1165665600, 1165669200, 1165672800, 1165676400, 1165680000, 
    1165683600, 1165687200, 1165690800, 1165694400, 1165698000, 1165701600, 
    1165705200, 1165708800, 1165712400, 1165716000, 1165719600, 1165723200, 
    1165726800, 1165730400, 1165734000, 1165737600, 1165741200, 1165744800, 
    1165748400, 1165752000, 1165755600, 1165759200, 1165762800, 1165766400, 
    1165770000, 1165773600, 1165777200, 1165780800, 1165784400, 1165788000, 
    1165791600, 1165795200, 1165798800, 1165802400, 1165806000, 1165809600, 
    1165813200, 1165816800, 1165820400, 1165824000, 1165827600, 1165831200, 
    1165834800, 1165838400, 1165842000, 1165845600, 1165849200, 1165852800, 
    1165856400, 1165860000, 1165863600, 1165867200, 1165870800, 1165874400, 
    1165878000, 1165881600, 1165885200, 1165888800, 1165892400, 1165896000, 
    1165899600, 1165903200, 1165906800, 1165910400, 1165914000, 1165917600, 
    1165921200, 1165924800, 1165928400, 1165932000, 1165935600, 1165939200, 
    1165942800, 1165946400, 1165950000, 1165953600, 1165957200, 1165960800, 
    1165964400, 1165968000, 1165971600, 1165975200, 1165978800, 1165982400, 
    1165986000, 1165989600, 1165993200, 1165996800, 1166000400, 1166004000, 
    1166007600, 1166011200, 1166014800, 1166018400, 1166022000, 1166025600, 
    1166029200, 1166032800, 1166036400, 1166040000, 1166043600, 1166047200, 
    1166050800, 1166054400, 1166058000, 1166061600, 1166065200, 1166068800, 
    1166072400, 1166076000, 1166079600, 1166083200, 1166086800, 1166090400, 
    1166094000, 1166097600, 1166101200, 1166104800, 1166108400, 1166112000, 
    1166115600, 1166119200, 1166122800, 1166126400, 1166130000, 1166133600, 
    1166137200, 1166140800, 1166144400, 1166148000, 1166151600, 1166155200, 
    1166158800, 1166162400, 1166166000, 1166169600, 1166173200, 1166176800, 
    1166180400, 1166184000, 1166187600, 1166191200, 1166194800, 1166198400, 
    1166202000, 1166205600, 1166209200, 1166212800, 1166216400, 1166220000, 
    1166223600, 1166227200, 1166230800, 1166234400, 1166238000, 1166241600, 
    1166245200, 1166248800, 1166252400, 1166256000, 1166259600, 1166263200, 
    1166266800, 1166270400, 1166274000, 1166277600, 1166281200, 1166284800, 
    1166288400, 1166292000, 1166295600, 1166299200, 1166302800, 1166306400, 
    1166310000, 1166313600, 1166317200, 1166320800, 1166324400, 1166328000, 
    1166331600, 1166335200, 1166338800, 1166342400, 1166346000, 1166349600, 
    1166353200, 1166356800, 1166360400, 1166364000, 1166367600, 1166371200, 
    1166374800, 1166378400, 1166382000, 1166385600, 1166389200, 1166392800, 
    1166396400, 1166400000, 1166403600, 1166407200, 1166410800, 1166414400, 
    1166418000, 1166421600, 1166425200, 1166428800, 1166432400, 1166436000, 
    1166439600, 1166443200, 1166446800, 1166450400, 1166454000, 1166457600, 
    1166461200, 1166464800, 1166468400, 1166472000, 1166475600, 1166479200, 
    1166482800, 1166486400, 1166490000, 1166493600, 1166497200, 1166500800, 
    1166504400, 1166508000, 1166511600, 1166515200, 1166518800, 1166522400, 
    1166526000, 1166529600, 1166533200, 1166536800, 1166540400, 1166544000, 
    1166547600, 1166551200, 1166554800, 1166558400, 1166562000, 1166565600, 
    1166569200, 1166572800, 1166576400, 1166580000, 1166583600, 1166587200, 
    1166590800, 1166594400, 1166598000, 1166601600, 1166605200, 1166608800, 
    1166612400, 1166616000, 1166619600, 1166623200, 1166626800, 1166630400, 
    1166634000, 1166637600, 1166641200, 1166644800, 1166648400, 1166652000, 
    1166655600, 1166659200, 1166662800, 1166666400, 1166670000, 1166673600, 
    1166677200, 1166680800, 1166684400, 1166688000, 1166691600, 1166695200, 
    1166698800, 1166702400, 1166706000, 1166709600, 1166713200, 1166716800, 
    1166720400, 1166724000, 1166727600, 1166731200, 1166734800, 1166738400, 
    1166742000, 1166745600, 1166749200, 1166752800, 1166756400, 1166760000, 
    1166763600, 1166767200, 1166770800, 1166774400, 1166778000, 1166781600, 
    1166785200, 1166788800, 1166792400, 1166796000, 1166799600, 1166803200, 
    1166806800, 1166810400, 1166814000, 1166817600, 1166821200, 1166824800, 
    1166828400, 1166832000, 1166835600, 1166839200, 1166842800, 1166846400, 
    1166850000, 1166853600, 1166857200, 1166860800, 1166864400, 1166868000, 
    1166871600, 1166875200, 1166878800, 1166882400, 1166886000, 1166889600, 
    1166893200, 1166896800, 1166900400, 1166904000, 1166907600, 1166911200, 
    1166914800, 1166918400, 1166922000, 1166925600, 1166929200, 1166932800, 
    1166936400, 1166940000, 1166943600, 1166947200, 1166950800, 1166954400, 
    1166958000, 1166961600, 1166965200, 1166968800, 1166972400, 1166976000, 
    1166979600, 1166983200, 1166986800, 1166990400, 1166994000, 1166997600, 
    1167001200, 1167004800, 1167008400, 1167012000, 1167015600, 1167019200, 
    1167022800, 1167026400, 1167030000, 1167033600, 1167037200, 1167040800, 
    1167044400, 1167048000, 1167051600, 1167055200, 1167058800, 1167062400, 
    1167066000, 1167069600, 1167073200, 1167076800, 1167080400, 1167084000, 
    1167087600, 1167091200, 1167094800, 1167098400, 1167102000, 1167105600, 
    1167109200, 1167112800, 1167116400, 1167120000, 1167123600, 1167127200, 
    1167130800, 1167134400, 1167138000, 1167141600, 1167145200, 1167148800, 
    1167152400, 1167156000, 1167159600, 1167163200, 1167166800, 1167170400, 
    1167174000, 1167177600, 1167181200, 1167184800, 1167188400, 1167192000, 
    1167195600, 1167199200, 1167202800, 1167206400, 1167210000, 1167213600, 
    1167217200, 1167220800, 1167224400, 1167228000, 1167231600, 1167235200, 
    1167238800, 1167242400, 1167246000, 1167249600, 1167253200, 1167256800, 
    1167260400, 1167264000, 1167267600, 1167271200, 1167274800, 1167278400, 
    1167282000, 1167285600, 1167289200, 1167292800, 1167296400, 1167300000, 
    1167303600, 1167307200, 1167310800, 1167314400, 1167318000, 1167321600, 
    1167325200, 1167328800, 1167332400, 1167336000, 1167339600, 1167343200, 
    1167346800, 1167350400, 1167354000, 1167357600, 1167361200, 1167364800, 
    1167368400, 1167372000, 1167375600, 1167379200, 1167382800, 1167386400, 
    1167390000, 1167393600, 1167397200, 1167400800, 1167404400, 1167408000, 
    1167411600, 1167415200, 1167418800, 1167422400, 1167426000, 1167429600, 
    1167433200, 1167436800, 1167440400, 1167444000, 1167447600, 1167451200, 
    1167454800, 1167458400, 1167462000, 1167465600, 1167469200, 1167472800, 
    1167476400, 1167480000, 1167483600, 1167487200, 1167490800, 1167494400, 
    1167498000, 1167501600, 1167505200, 1167508800, 1167512400, 1167516000, 
    1167519600, 1167523200, 1167526800, 1167530400, 1167534000, 1167537600, 
    1167541200, 1167544800, 1167548400, 1167552000, 1167555600, 1167559200, 
    1167562800, 1167566400, 1167570000, 1167573600, 1167577200, 1167580800, 
    1167584400, 1167588000, 1167591600, 1167595200, 1167598800, 1167602400, 
    1167606000, 1167609600, 1167613200, 1167616800, 1167620400, 1167624000, 
    1167627600, 1167631200, 1167634800, 1167638400, 1167642000, 1167645600, 
    1167649200, 1167652800, 1167656400, 1167660000, 1167663600, 1167667200, 
    1167670800, 1167674400, 1167678000, 1167681600, 1167685200, 1167688800, 
    1167692400, 1167696000, 1167699600, 1167703200, 1167706800, 1167710400, 
    1167714000, 1167717600, 1167721200, 1167724800, 1167728400, 1167732000, 
    1167735600, 1167739200, 1167742800, 1167746400, 1167750000, 1167753600, 
    1167757200, 1167760800, 1167764400, 1167768000, 1167771600, 1167775200, 
    1167778800, 1167782400, 1167786000, 1167789600, 1167793200, 1167796800, 
    1167800400, 1167804000, 1167807600, 1167811200, 1167814800, 1167818400, 
    1167822000, 1167825600, 1167829200, 1167832800, 1167836400, 1167840000, 
    1167843600, 1167847200, 1167850800, 1167854400, 1167858000, 1167861600, 
    1167865200, 1167868800, 1167872400, 1167876000, 1167879600, 1167883200, 
    1167886800, 1167890400, 1167894000, 1167897600, 1167901200, 1167904800, 
    1167908400, 1167912000, 1167915600, 1167919200, 1167922800, 1167926400, 
    1167930000, 1167933600, 1167937200, 1167940800, 1167944400, 1167948000, 
    1167951600, 1167955200, 1167958800, 1167962400, 1167966000, 1167969600, 
    1167973200, 1167976800, 1167980400, 1167984000, 1167987600, 1167991200, 
    1167994800, 1167998400, 1168002000, 1168005600, 1168009200, 1168012800, 
    1168016400, 1168020000, 1168023600, 1168027200, 1168030800, 1168034400, 
    1168038000, 1168041600, 1168045200, 1168048800, 1168052400, 1168056000, 
    1168059600, 1168063200, 1168066800, 1168070400, 1168074000, 1168077600, 
    1168081200, 1168084800, 1168088400, 1168092000, 1168095600, 1168099200, 
    1168102800, 1168106400, 1168110000, 1168113600, 1168117200, 1168120800, 
    1168124400, 1168128000, 1168131600, 1168135200, 1168138800, 1168142400, 
    1168146000, 1168149600, 1168153200, 1168156800, 1168160400, 1168164000, 
    1168167600, 1168171200, 1168174800, 1168178400, 1168182000, 1168185600, 
    1168189200, 1168192800, 1168196400, 1168200000, 1168203600, 1168207200, 
    1168210800, 1168214400, 1168218000, 1168221600, 1168225200, 1168228800, 
    1168232400, 1168236000, 1168239600, 1168243200, 1168246800, 1168250400, 
    1168254000, 1168257600, 1168261200, 1168264800, 1168268400, 1168272000, 
    1168275600, 1168279200, 1168282800, 1168286400, 1168290000, 1168293600, 
    1168297200, 1168300800, 1168304400, 1168308000, 1168311600, 1168315200, 
    1168318800, 1168322400, 1168326000, 1168329600, 1168333200, 1168336800, 
    1168340400, 1168344000, 1168347600, 1168351200, 1168354800, 1168358400, 
    1168362000, 1168365600, 1168369200, 1168372800, 1168376400, 1168380000, 
    1168383600, 1168387200, 1168390800, 1168394400, 1168398000, 1168401600, 
    1168405200, 1168408800, 1168412400, 1168416000, 1168419600, 1168423200, 
    1168426800, 1168430400, 1168434000, 1168437600, 1168441200, 1168444800, 
    1168448400, 1168452000, 1168455600, 1168459200, 1168462800, 1168466400, 
    1168470000, 1168473600, 1168477200, 1168480800, 1168484400, 1168488000, 
    1168491600, 1168495200, 1168498800, 1168502400, 1168506000, 1168509600, 
    1168513200, 1168516800, 1168520400, 1168524000, 1168527600, 1168531200, 
    1168534800, 1168538400, 1168542000, 1168545600, 1168549200, 1168552800, 
    1168556400, 1168560000, 1168563600, 1168567200, 1168570800, 1168574400, 
    1168578000, 1168581600, 1168585200, 1168588800, 1168592400, 1168596000, 
    1168599600, 1168603200, 1168606800, 1168610400, 1168614000, 1168617600, 
    1168621200, 1168624800, 1168628400, 1168632000, 1168635600, 1168639200, 
    1168642800, 1168646400, 1168650000, 1168653600, 1168657200, 1168660800, 
    1168664400, 1168668000, 1168671600, 1168675200, 1168678800, 1168682400, 
    1168686000, 1168689600, 1168693200, 1168696800, 1168700400, 1168704000, 
    1168707600, 1168711200, 1168714800, 1168718400, 1168722000, 1168725600, 
    1168729200, 1168732800, 1168736400, 1168740000, 1168743600, 1168747200, 
    1168750800, 1168754400, 1168758000, 1168761600, 1168765200, 1168768800, 
    1168772400, 1168776000, 1168779600, 1168783200, 1168786800, 1168790400, 
    1168794000, 1168797600, 1168801200, 1168804800, 1168808400, 1168812000, 
    1168815600, 1168819200, 1168822800, 1168826400, 1168830000, 1168833600, 
    1168837200, 1168840800, 1168844400, 1168848000, 1168851600, 1168855200, 
    1168858800, 1168862400, 1168866000, 1168869600, 1168873200, 1168876800, 
    1168880400, 1168884000, 1168887600, 1168891200, 1168894800, 1168898400, 
    1168902000, 1168905600, 1168909200, 1168912800, 1168916400, 1168920000, 
    1168923600, 1168927200, 1168930800, 1168934400, 1168938000, 1168941600, 
    1168945200, 1168948800, 1168952400, 1168956000, 1168959600, 1168963200, 
    1168966800, 1168970400, 1168974000, 1168977600, 1168981200, 1168984800, 
    1168988400, 1168992000, 1168995600, 1168999200, 1169002800, 1169006400, 
    1169010000, 1169013600, 1169017200, 1169020800, 1169024400, 1169028000, 
    1169031600, 1169035200, 1169038800, 1169042400, 1169046000, 1169049600, 
    1169053200, 1169056800, 1169060400, 1169064000, 1169067600, 1169071200, 
    1169074800, 1169078400, 1169082000, 1169085600, 1169089200, 1169092800, 
    1169096400, 1169100000, 1169103600, 1169107200, 1169110800, 1169114400, 
    1169118000, 1169121600, 1169125200, 1169128800, 1169132400, 1169136000, 
    1169139600, 1169143200, 1169146800, 1169150400, 1169154000, 1169157600, 
    1169161200, 1169164800, 1169168400, 1169172000, 1169175600, 1169179200, 
    1169182800, 1169186400, 1169190000, 1169193600, 1169197200, 1169200800, 
    1169204400, 1169208000, 1169211600, 1169215200, 1169218800, 1169222400, 
    1169226000, 1169229600, 1169233200, 1169236800, 1169240400, 1169244000, 
    1169247600, 1169251200, 1169254800, 1169258400, 1169262000, 1169265600, 
    1169269200, 1169272800, 1169276400, 1169280000, 1169283600, 1169287200, 
    1169290800, 1169294400, 1169298000, 1169301600, 1169305200, 1169308800, 
    1169312400, 1169316000, 1169319600, 1169323200, 1169326800, 1169330400, 
    1169334000, 1169337600, 1169341200, 1169344800, 1169348400, 1169352000, 
    1169355600, 1169359200, 1169362800, 1169366400, 1169370000, 1169373600, 
    1169377200, 1169380800, 1169384400, 1169388000, 1169391600, 1169395200, 
    1169398800, 1169402400, 1169406000, 1169409600, 1169413200, 1169416800, 
    1169420400, 1169424000, 1169427600, 1169431200, 1169434800, 1169438400, 
    1169442000, 1169445600, 1169449200, 1169452800, 1169456400, 1169460000, 
    1169463600, 1169467200, 1169470800, 1169474400, 1169478000, 1169481600, 
    1169485200, 1169488800, 1169492400, 1169496000, 1169499600, 1169503200, 
    1169506800, 1169510400, 1169514000, 1169517600, 1169521200, 1169524800, 
    1169528400, 1169532000, 1169535600, 1169539200, 1169542800, 1169546400, 
    1169550000, 1169553600, 1169557200, 1169560800, 1169564400, 1169568000, 
    1169571600, 1169575200, 1169578800, 1169582400, 1169586000, 1169589600, 
    1169593200, 1169596800, 1169600400, 1169604000, 1169607600, 1169611200, 
    1169614800, 1169618400, 1169622000, 1169625600, 1169629200, 1169632800, 
    1169636400, 1169640000, 1169643600, 1169647200, 1169650800, 1169654400, 
    1169658000, 1169661600, 1169665200, 1169668800, 1169672400, 1169676000, 
    1169679600, 1169683200, 1169686800, 1169690400, 1169694000, 1169697600, 
    1169701200, 1169704800, 1169708400, 1169712000, 1169715600, 1169719200, 
    1169722800, 1169726400, 1169730000, 1169733600, 1169737200, 1169740800, 
    1169744400, 1169748000, 1169751600, 1169755200, 1169758800, 1169762400, 
    1169766000, 1169769600, 1169773200, 1169776800, 1169780400, 1169784000, 
    1169787600, 1169791200, 1169794800, 1169798400, 1169802000, 1169805600, 
    1169809200, 1169812800, 1169816400, 1169820000, 1169823600, 1169827200, 
    1169830800, 1169834400, 1169838000, 1169841600, 1169845200, 1169848800, 
    1169852400, 1169856000, 1169859600, 1169863200, 1169866800, 1169870400, 
    1169874000, 1169877600, 1169881200, 1169884800, 1169888400, 1169892000, 
    1169895600, 1169899200, 1169902800, 1169906400, 1169910000, 1169913600, 
    1169917200, 1169920800, 1169924400, 1169928000, 1169931600, 1169935200, 
    1169938800, 1169942400, 1169946000, 1169949600, 1169953200, 1169956800, 
    1169960400, 1169964000, 1169967600, 1169971200, 1169974800, 1169978400, 
    1169982000, 1169985600, 1169989200, 1169992800, 1169996400, 1170000000, 
    1170003600, 1170007200, 1170010800, 1170014400, 1170018000, 1170021600, 
    1170025200, 1170028800, 1170032400, 1170036000, 1170039600, 1170043200, 
    1170046800, 1170050400, 1170054000, 1170057600, 1170061200, 1170064800, 
    1170068400, 1170072000, 1170075600, 1170079200, 1170082800, 1170086400, 
    1170090000, 1170093600, 1170097200, 1170100800, 1170104400, 1170108000, 
    1170111600, 1170115200, 1170118800, 1170122400, 1170126000, 1170129600, 
    1170133200, 1170136800, 1170140400, 1170144000, 1170147600, 1170151200, 
    1170154800, 1170158400, 1170162000, 1170165600, 1170169200, 1170172800, 
    1170176400, 1170180000, 1170183600, 1170187200, 1170190800, 1170194400, 
    1170198000, 1170201600, 1170205200, 1170208800, 1170212400, 1170216000, 
    1170219600, 1170223200, 1170226800, 1170230400, 1170234000, 1170237600, 
    1170241200, 1170244800, 1170248400, 1170252000, 1170255600, 1170259200, 
    1170262800, 1170266400, 1170270000, 1170273600, 1170277200, 1170280800, 
    1170284400, 1170288000, 1170291600, 1170295200, 1170298800, 1170302400, 
    1170306000, 1170309600, 1170313200, 1170316800, 1170320400, 1170324000, 
    1170327600, 1170331200, 1170334800, 1170338400, 1170342000, 1170345600, 
    1170349200, 1170352800, 1170356400, 1170360000, 1170363600, 1170367200, 
    1170370800, 1170374400, 1170378000, 1170381600, 1170385200, 1170388800, 
    1170392400, 1170396000, 1170399600, 1170403200, 1170406800, 1170410400, 
    1170414000, 1170417600, 1170421200, 1170424800, 1170428400, 1170432000, 
    1170435600, 1170439200, 1170442800, 1170446400, 1170450000, 1170453600, 
    1170457200, 1170460800, 1170464400, 1170468000, 1170471600, 1170475200, 
    1170478800, 1170482400, 1170486000, 1170489600, 1170493200, 1170496800, 
    1170500400, 1170504000, 1170507600, 1170511200, 1170514800, 1170518400, 
    1170522000, 1170525600, 1170529200, 1170532800, 1170536400, 1170540000, 
    1170543600, 1170547200, 1170550800, 1170554400, 1170558000, 1170561600, 
    1170565200, 1170568800, 1170572400, 1170576000, 1170579600, 1170583200, 
    1170586800, 1170590400, 1170594000, 1170597600, 1170601200, 1170604800, 
    1170608400, 1170612000, 1170615600, 1170619200, 1170622800, 1170626400, 
    1170630000, 1170633600, 1170637200, 1170640800, 1170644400, 1170648000, 
    1170651600, 1170655200, 1170658800, 1170662400, 1170666000, 1170669600, 
    1170673200, 1170676800, 1170680400, 1170684000, 1170687600, 1170691200, 
    1170694800, 1170698400, 1170702000, 1170705600, 1170709200, 1170712800, 
    1170716400, 1170720000, 1170723600, 1170727200, 1170730800, 1170734400, 
    1170738000, 1170741600, 1170745200, 1170748800, 1170752400, 1170756000, 
    1170759600, 1170763200, 1170766800, 1170770400, 1170774000, 1170777600, 
    1170781200, 1170784800, 1170788400, 1170792000, 1170795600, 1170799200, 
    1170802800, 1170806400, 1170810000, 1170813600, 1170817200, 1170820800, 
    1170824400, 1170828000, 1170831600, 1170835200, 1170838800, 1170842400, 
    1170846000, 1170849600, 1170853200, 1170856800, 1170860400, 1170864000, 
    1170867600, 1170871200, 1170874800, 1170878400, 1170882000, 1170885600, 
    1170889200, 1170892800, 1170896400, 1170900000, 1170903600, 1170907200, 
    1170910800, 1170914400, 1170918000, 1170921600, 1170925200, 1170928800, 
    1170932400, 1170936000, 1170939600, 1170943200, 1170946800, 1170950400, 
    1170954000, 1170957600, 1170961200, 1170964800, 1170968400, 1170972000, 
    1170975600, 1170979200, 1170982800, 1170986400, 1170990000, 1170993600, 
    1170997200, 1171000800, 1171004400, 1171008000, 1171011600, 1171015200, 
    1171018800, 1171022400, 1171026000, 1171029600, 1171033200, 1171036800, 
    1171040400, 1171044000, 1171047600, 1171051200, 1171054800, 1171058400, 
    1171062000, 1171065600, 1171069200, 1171072800, 1171076400, 1171080000, 
    1171083600, 1171087200, 1171090800, 1171094400, 1171098000, 1171101600, 
    1171105200, 1171108800, 1171112400, 1171116000, 1171119600, 1171123200, 
    1171126800, 1171130400, 1171134000, 1171137600, 1171141200, 1171144800, 
    1171148400, 1171152000, 1171155600, 1171159200, 1171162800, 1171166400, 
    1171170000, 1171173600, 1171177200, 1171180800, 1171184400, 1171188000, 
    1171191600, 1171195200, 1171198800, 1171202400, 1171206000, 1171209600, 
    1171213200, 1171216800, 1171220400, 1171224000, 1171227600, 1171231200, 
    1171234800, 1171238400, 1171242000, 1171245600, 1171249200, 1171252800, 
    1171256400, 1171260000, 1171263600, 1171267200, 1171270800, 1171274400, 
    1171278000, 1171281600, 1171285200, 1171288800, 1171292400, 1171296000, 
    1171299600, 1171303200, 1171306800, 1171310400, 1171314000, 1171317600, 
    1171321200, 1171324800, 1171328400, 1171332000, 1171335600, 1171339200, 
    1171342800, 1171346400, 1171350000, 1171353600, 1171357200, 1171360800, 
    1171364400, 1171368000, 1171371600, 1171375200, 1171378800, 1171382400, 
    1171386000, 1171389600, 1171393200, 1171396800, 1171400400, 1171404000, 
    1171407600, 1171411200, 1171414800, 1171418400, 1171422000, 1171425600, 
    1171429200, 1171432800, 1171436400, 1171440000, 1171443600, 1171447200, 
    1171450800, 1171454400, 1171458000, 1171461600, 1171465200, 1171468800, 
    1171472400, 1171476000, 1171479600, 1171483200, 1171486800, 1171490400, 
    1171494000, 1171497600, 1171501200, 1171504800, 1171508400, 1171512000, 
    1171515600, 1171519200, 1171522800, 1171526400, 1171530000, 1171533600, 
    1171537200, 1171540800, 1171544400, 1171548000, 1171551600, 1171555200, 
    1171558800, 1171562400, 1171566000, 1171569600, 1171573200, 1171576800, 
    1171580400, 1171584000, 1171587600, 1171591200, 1171594800, 1171598400, 
    1171602000, 1171605600, 1171609200, 1171612800, 1171616400, 1171620000, 
    1171623600, 1171627200, 1171630800, 1171634400, 1171638000, 1171641600, 
    1171645200, 1171648800, 1171652400, 1171656000, 1171659600, 1171663200, 
    1171666800, 1171670400, 1171674000, 1171677600, 1171681200, 1171684800, 
    1171688400, 1171692000, 1171695600, 1171699200, 1171702800, 1171706400, 
    1171710000, 1171713600, 1171717200, 1171720800, 1171724400, 1171728000, 
    1171731600, 1171735200, 1171738800, 1171742400, 1171746000, 1171749600, 
    1171753200, 1171756800, 1171760400, 1171764000, 1171767600, 1171771200, 
    1171774800, 1171778400, 1171782000, 1171785600, 1171789200, 1171792800, 
    1171796400, 1171800000, 1171803600, 1171807200, 1171810800, 1171814400, 
    1171818000, 1171821600, 1171825200, 1171828800, 1171832400, 1171836000, 
    1171839600, 1171843200, 1171846800, 1171850400, 1171854000, 1171857600, 
    1171861200, 1171864800, 1171868400, 1171872000, 1171875600, 1171879200, 
    1171882800, 1171886400, 1171890000, 1171893600, 1171897200, 1171900800, 
    1171904400, 1171908000, 1171911600, 1171915200, 1171918800, 1171922400, 
    1171926000, 1171929600, 1171933200, 1171936800, 1171940400, 1171944000, 
    1171947600, 1171951200, 1171954800, 1171958400, 1171962000, 1171965600, 
    1171969200, 1171972800, 1171976400, 1171980000, 1171983600, 1171987200, 
    1171990800, 1171994400, 1171998000, 1172001600, 1172005200, 1172008800, 
    1172012400, 1172016000, 1172019600, 1172023200, 1172026800, 1172030400, 
    1172034000, 1172037600, 1172041200, 1172044800, 1172048400, 1172052000, 
    1172055600, 1172059200, 1172062800, 1172066400, 1172070000, 1172073600, 
    1172077200, 1172080800, 1172084400, 1172088000, 1172091600, 1172095200, 
    1172098800, 1172102400, 1172106000, 1172109600, 1172113200, 1172116800, 
    1172120400, 1172124000, 1172127600, 1172131200, 1172134800, 1172138400, 
    1172142000, 1172145600, 1172149200, 1172152800, 1172156400, 1172160000, 
    1172163600, 1172167200, 1172170800, 1172174400, 1172178000, 1172181600, 
    1172185200, 1172188800, 1172192400, 1172196000, 1172199600, 1172203200, 
    1172206800, 1172210400, 1172214000, 1172217600, 1172221200, 1172224800, 
    1172228400, 1172232000, 1172235600, 1172239200, 1172242800, 1172246400, 
    1172250000, 1172253600, 1172257200, 1172260800, 1172264400, 1172268000, 
    1172271600, 1172275200, 1172278800, 1172282400, 1172286000, 1172289600, 
    1172293200, 1172296800, 1172300400, 1172304000, 1172307600, 1172311200, 
    1172314800, 1172318400, 1172322000, 1172325600, 1172329200, 1172332800, 
    1172336400, 1172340000, 1172343600, 1172347200, 1172350800, 1172354400, 
    1172358000, 1172361600, 1172365200, 1172368800, 1172372400, 1172376000, 
    1172379600, 1172383200, 1172386800, 1172390400, 1172394000, 1172397600, 
    1172401200, 1172404800, 1172408400, 1172412000, 1172415600, 1172419200, 
    1172422800, 1172426400, 1172430000, 1172433600, 1172437200, 1172440800, 
    1172444400, 1172448000, 1172451600, 1172455200, 1172458800, 1172462400, 
    1172466000, 1172469600, 1172473200, 1172476800, 1172480400, 1172484000, 
    1172487600, 1172491200, 1172494800, 1172498400, 1172502000, 1172505600, 
    1172509200, 1172512800, 1172516400, 1172520000, 1172523600, 1172527200, 
    1172530800, 1172534400, 1172538000, 1172541600, 1172545200, 1172548800, 
    1172552400, 1172556000, 1172559600, 1172563200, 1172566800, 1172570400, 
    1172574000, 1172577600, 1172581200, 1172584800, 1172588400, 1172592000, 
    1172595600, 1172599200, 1172602800, 1172606400, 1172610000, 1172613600, 
    1172617200, 1172620800, 1172624400, 1172628000, 1172631600, 1172635200, 
    1172638800, 1172642400, 1172646000, 1172649600, 1172653200, 1172656800, 
    1172660400, 1172664000, 1172667600, 1172671200, 1172674800, 1172678400, 
    1172682000, 1172685600, 1172689200, 1172692800, 1172696400, 1172700000, 
    1172703600 ;

 Prec =
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.6, 0.8, 1.2},
  {0.8, 1, 1.4},
  {0.4, 0.8, 1.2},
  {0.4, 1, 1},
  {0.6, 0.8, 1.4},
  {0.4, 0.6, 1.2},
  {0, 0, 0.6},
  {0.4, 0, 0.2},
  {0.2, 0, 0.4},
  {0.8, 0.2, 0.4},
  {0.2, 0.2, 0.2},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.8, 0, 0.6},
  {0, 0.2, 0},
  {0, 0.6, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.8, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0.4, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 2.4, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 1, 0},
  {0.2, 1.2, 0},
  {0.6, 2.4, 0.8},
  {0, 0.4, 1.4},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 2.6, 0},
  {0, 0.4, 0},
  {0, 0.2, 0.4},
  {0.2, 0, 1},
  {0.4, 0, 0},
  {0.4, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0.2},
  {6.2, 0, 0.6},
  {0, 0, 0.2},
  {0, 0, 0},
  {0.4, 0, 0},
  {0, 0, 0.2},
  {0, 0.6, 0},
  {0, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0.2},
  {2, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0.2, 0},
  {0, 0.2, 0.2},
  {0, 0, 0.4},
  {1.4, 0.2, 1.4},
  {2, 0.4, 2},
  {3, 2.2, 4},
  {2.6, 3.4, 4.4},
  {3.2, 2.4, 4.4},
  {4, 3.2, 6},
  {3.2, 3.6, 6.2},
  {2.8, 2.8, 5},
  {2.2, 1.8, 1.4},
  {2.4, 2.6, 1.2},
  {2.2, 0.4, 0.6},
  {1, 0.6, 0.2},
  {0.4, 0.4, 0.6},
  {0, 1, 0.2},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.8, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.6, 0, 0},
  {0.4, 0, 0},
  {0.8, 0, 0},
  {1.6, 0, 0},
  {1.4, 0, 0},
  {0.8, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.6, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1, 0, 0},
  {0.4, 0, 0.6},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {3.6, 0, 0.2},
  {5.2, 4.4, 5.8},
  {4.6, 2.4, 3.8},
  {5, 3.6, 3.6},
  {4.2, 2.8, 2.8},
  {4.8, 3, 4.8},
  {0.8, 4, 2.2},
  {0, 1.6, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.4, 0},
  {0, 0.6, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.6, 0, 0},
  {2.2, 0, 0.2},
  {1, 0, 1},
  {1, 0.8, 0.2},
  {1, 1.6, 0.6},
  {0.4, 2.2, 0.2},
  {0.4, 0, 0.2},
  {0.8, 0.4, 0},
  {2, 0.2, 0.2},
  {0, 0.6, 0},
  {0.2, 0.6, 0.6},
  {0, 0.8, 0.2},
  {0, 1.4, 0.4},
  {0, 3, 0.2},
  {0, 3.2, 0.2},
  {0, 1.2, 1.6},
  {0, 0.4, 1},
  {0, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0.6, 0, 0},
  {0.8, 0, 0},
  {0, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1, 0.4, 0.2},
  {1.2, 1.6, 2.4},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1, 0, 0.4},
  {1.4, 0.8, 1.6},
  {2.2, 1, 2.2},
  {1.6, 2.2, 3.2},
  {0.8, 1.8, 1},
  {0.8, 1.6, 1.8},
  {0.2, 0.4, 0.4},
  {0, 0.2, 0.2},
  {0, 0, 0},
  {0.4, 0, 0},
  {0.8, 0.2, 0.4},
  {2.6, 0.2, 0},
  {0.6, 0, 0},
  {0.2, 0, 0},
  {0.2, 0.2, 0},
  {0, 1.8, 1.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0.8, 0.2, 1},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {_, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1.2, 0.2, 0},
  {1.4, 8.6, 5.6},
  {0, 6.2, 0.2},
  {0, 0.6, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.6, 0, 0},
  {1, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {1, 0, 0.2},
  {1, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, _},
  {0, 0, _},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 1.6, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {3.2, 0, 0},
  {1.6, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0.2, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {2.4, 0, 0},
  {1.6, 0.4, 0},
  {1.6, 0.4, 0.8},
  {3.2, 0.2, 0.6},
  {6.6, 0.4, 2},
  {0.6, 0.2, 1.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1.4, 0, 0},
  {0.8, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 1.4},
  {0.8, 0.4, 3.8},
  {2, 3, 1},
  {1.8, 2.8, 0.2},
  {0, 3.4, 0.2},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.4, 0},
  {0, 1.8, 0.2},
  {0, 0, 0},
  {0.6, 0, 0},
  {5, 0, 0.8},
  {1.6, 0.8, 5},
  {2.2, 2, 2.4},
  {1.8, 0.6, 2.2},
  {3, 2.6, 2.8},
  {2.4, 4.2, 5},
  {1.6, 3, 4},
  {0.8, 3, 1.4},
  {3.2, 5, 2.4},
  {0.8, 5.4, 1.8},
  {5.8, 3.2, 1.6},
  {6.2, 3.8, 7.6},
  {1.8, 5.6, 5.6},
  {0.4, 5, 5},
  {1.2, 4, 3.8},
  {0.8, 1.4, 2},
  {1, 0, 0.8},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.6},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0.6, 0.4, 1.6},
  {1.2, 1.6, 2},
  {0, 0.2, 0.2},
  {0, 0.6, 0},
  {0.6, 2.4, 1.4},
  {0.2, 0, 1.8},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 1, 0},
  {0, 3, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0.4, 5.8},
  {0, 0, 7},
  {0, 0, 1.6},
  {0, 0.2, 0},
  {0, 1.8, 0},
  {0, 0, 0},
  {0, 1.2, 0},
  {0, 0.2, 0},
  {0.4, 0, 0},
  {0.4, 0, 0},
  {1, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.4, 0},
  {0, 0.8, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 6.6},
  {4.2, 0, 2},
  {1.6, 0, 0.4},
  {0.2, 0, 0.2},
  {0, 0, 0.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, 0.8},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 3},
  {0.2, 0, 4.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {5.6, 0.4, 1.2},
  {0, 0, 4.4},
  {0.2, 0.4, 0.2},
  {1.6, 0.4, 0.8},
  {0.6, 0.4, 1.6},
  {0, 0.4, 1},
  {0.2, 0, 0},
  {0.2, 0, 0.6},
  {0, 0.4, 0},
  {0.2, 0.8, 1},
  {0.2, 2, 0.8},
  {0, 2.6, 0.6},
  {0, 1.6, 0.2},
  {0, 2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1.2, 0, 0},
  {0, 17.4, 0.8},
  {0, 0.4, 1},
  {0, 0.2, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.8},
  {0, 0, 2.4},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 1, 4.6},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {2.4, 0, 0},
  {0.6, 0, 0},
  {1.2, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {9.8, 0, 0.2},
  {6.6, 0, 1.6},
  {8.8, 0, 0.2},
  {1, 0, 0},
  {0.6, 0, 2.2},
  {1, 0, 1.6},
  {0, 0, 1},
  {0, 2.6, 0.2},
  {4, 11.6, 4.4},
  {6.2, 4.8, 14.2},
  {0, 0.2, 0},
  {1.2, 1.4, 0.6},
  {1, 0, 0.2},
  {4.4, 0, 0.2},
  {4.2, 3, 4.6},
  {0, 0.6, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.8, 6.2, 0.2},
  {6.8, 1.4, 3.2},
  {0, 0.2, 2.4},
  {0.2, 0, 0.8},
  {0, 0, 0},
  {0.8, 1.6, 1},
  {0.4, 0.8, 0.6},
  {0, 0.2, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.4, 0},
  {1, 0.2, 1.4},
  {0.4, 0.6, 0.6},
  {3, 0.4, 1.8},
  {0.4, 3.8, 3.4},
  {0.2, 0.6, 0.6},
  {0, 0, 0},
  {0, 0, 0},
  {1.4, 0, 1.2},
  {1.4, 1.6, 2.4},
  {0.4, 3.6, 0.4},
  {5.6, 1, 2.6},
  {2.4, 1.2, 2.2},
  {0.6, 0.4, 1.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1.2, 0, 0.4},
  {0.2, 0.8, 6.6},
  {0, 1.4, 2.2},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0.4, 0.6, 0},
  {1, 0, 0},
  {4.4, 0, 0},
  {1, 0, 0},
  {1, 4.6, 1.2},
  {1.4, 6.2, 4.4},
  {13.2, 7.6, 7.2},
  {5.6, 3.4, 4.2},
  {0.2, 3.4, 1.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0.6, 0},
  {0.2, 0.4, 0},
  {0.2, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 1.4, 0},
  {0, 0.4, 0.2},
  {0.2, 0, 0.6},
  {0.2, 0, 0.2},
  {0.6, 0, 0.2},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, _, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 1.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, _, 0},
  {0, 0.2, 0},
  {0, 8.4, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 1.2, 0},
  {10.6, 4.4, 7.8},
  {11.8, 1.4, 1.6},
  {0.2, 0.2, 0.8},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0.6},
  {14.8, 0, 1.8},
  {28, 0, 0},
  {3.8, 0, 0},
  {0.6, 0, 0},
  {0.6, 0.2, 0.4},
  {1.6, 3, 2.6},
  {1, 5, 1},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 7.4, 0},
  {0, 0.6, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1, 0, 0},
  {0, 0.8, 0},
  {0.2, 0.2, 0},
  {0, 0, 0},
  {0.4, 0.4, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0, 0, 0},
  {4.2, 3.4, 0.8},
  {3, 3.6, 6.8},
  {5.8, 4.4, 6},
  {2.6, 2.6, 2.4},
  {0, 7, 1.4},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.8, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 1.2, 0.2},
  {0, 0, 0.6},
  {0.2, 0, 0.4},
  {9.8, 0, 0},
  {1, 0, 0},
  {1.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, _},
  {0, 0, _},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 1.4, 10.2},
  {1.4, 3.2, 17.4},
  {0.4, 3.4, 0.8},
  {1, 0.4, 0.8},
  {0, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 1.4},
  {0.2, 0, 0},
  {0.4, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0.8, 0},
  {0, 0, 0.2},
  {0, 2, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {2, 0.2, 0.4},
  {0, 0, 0.4},
  {0.6, 0.6, 0.2},
  {3.2, 0, 5.4},
  {0.8, 0, 0.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {5.2, 0, 0.2},
  {4.6, 0.2, 0.8},
  {0.6, 1.4, 0},
  {0, 4, 0.4},
  {1.2, 5.8, 1.6},
  {0.8, 4, 0.2},
  {0, 1, 0},
  {1, 0, 0.8},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 1.2},
  {0, 0, 0},
  {0, 0.2, 0.2},
  {0.4, 0.8, 0.2},
  {2.4, 1.8, 1.6},
  {1.2, 1, 2.4},
  {0.8, 1, 2.8},
  {1.4, 1.4, 2},
  {2, 0.4, 1.8},
  {2.6, 0.2, 1.8},
  {2.2, 0, 1.2},
  {0.8, 0.6, 2.2},
  {0.2, 1.8, 1.4},
  {0.4, 0.6, 0.6},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0.2, 0, 0},
  {4.4, 0.6, 0},
  {1.6, 0.4, 1.8},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.6, 0},
  {0.8, 1, 0.4},
  {0.8, 0.2, 0.6},
  {0.4, 0.8, 0.2},
  {0, 0.4, 0.4},
  {0.2, 2.8, 1.2},
  {0.6, 1.4, 2.2},
  {0.6, 0, 0.6},
  {0, 0, 0},
  {0.4, 0.4, 0.2},
  {0.6, 1, 1.8},
  {1.2, 2, 2.6},
  {1, 0, 1.8},
  {0.4, 0.2, 1.2},
  {0.4, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0.4},
  {0, 0.4, 0.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1, 0, 0.4},
  {1.4, 0.4, 1.6},
  {0.6, 3.2, 1.4},
  {2.4, 9.6, 7.2},
  {0.6, 2.8, 4.4},
  {1, 0.8, 2.2},
  {0.2, 0, 1.4},
  {0, 0, 0.4},
  {0.8, 0, 0},
  {0.8, 0, 1},
  {1.6, 0, 0.2},
  {0.4, 0, 0.8},
  {0, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.4, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.4},
  {0, 0, 0},
  {0, 1.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0.2, 0, 0.4},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 1.6, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 1.6},
  {0.8, 0, 0.2},
  {0.6, 1.4, 10.8},
  {1.4, 3.6, 4.8},
  {0.2, 0.2, 0.8},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 1.6, 0},
  {0.8, 4.2, 0.8},
  {0.4, 2.6, 1},
  {1.2, 0.6, 1.6},
  {1.6, 4, 3.4},
  {0, 1.8, 4},
  {0, 0, 2.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 2.8, 0.4},
  {5.6, 3.8, 1.8},
  {5.2, 7.2, 7.4},
  {0.4, 2.4, 2.2},
  {0.2, 4, 1},
  {0, 0.2, 20},
  {0, 0, 1.6},
  {0.6, 0, 0.8},
  {0.2, 0.2, 5.8},
  {0.8, 0, 0.2},
  {0, 0.6, 0.2},
  {0, 0.6, 0},
  {1.8, 5.2, 0},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 3.6},
  {0, 8.8, 0.6},
  {0, 0.8, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0.2},
  {2.4, 0, 6.2},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.4},
  {0.2, 0, 0.2},
  {0.8, 8.4, 0.2},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0.8},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {3, 0, 1.6},
  {0, 1.8, 0.4},
  {5, 0.2, 1},
  {4.2, 0.8, 5.4},
  {2.6, 0.6, 1.2},
  {0.2, 0.6, 2},
  {0, 1.2, 1.4},
  {0, 0.2, 0.2},
  {0, 0.8, 0},
  {0, 0.4, 0},
  {0.4, 0.2, 0},
  {1, 1.8, 0},
  {1.2, 1, 0},
  {0.8, 1.2, 0.4},
  {0.4, 0.4, 0.2},
  {0.2, 0.4, 0},
  {0, 0, 0},
  {0.8, 0, 0},
  {0.8, 0.4, 0.6},
  {0.6, 0.6, 0.2},
  {0.2, 0.2, 0.2},
  {0.2, 0, 0.2},
  {0.2, 0.2, 0.2},
  {0.2, 0.4, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0.2, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0.2},
  {0, 0, 1},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 2},
  {0, 0.6, 0.2},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.2, 0, 0},
  {0, 4.4, 0},
  {0, 2.2, 0.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0.2, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0.4, 0.4},
  {0, 0.6, 0},
  {0, 0, 0.2},
  {0, 0.4, 0.6},
  {0.6, 0.2, 1.4},
  {0, 0.6, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0.4, 0, 1.4},
  {0.2, 0.4, 0.2},
  {1.4, 0.2, 0.6},
  {0.8, 1.4, 2.6},
  {0.4, 2, 2},
  {3, 1, 4.6},
  {0.8, 4, 4.8},
  {3.2, 5, 2.8},
  {0.8, 2.6, 3.2},
  {2.2, 1.2, 5},
  {4.2, 1.8, 4.8},
  {3.4, 3.2, 3.8},
  {6.2, 3.2, 8.2},
  {7, 3.2, 7.6},
  {2, 4.6, 3.6},
  {0, 2, 0.2},
  {0.4, 1.2, 0},
  {1.4, 3, 1.2},
  {0.4, 6.4, 0.8},
  {0.8, 3.2, 0.6},
  {0.4, 0.6, 0.8},
  {0.2, 0.2, 0},
  {0.2, 0, 1.6},
  {0.2, 0, 1},
  {0, 0, 0},
  {0, 0, 0},
  {0.8, 0.2, 0},
  {2.6, 2, 2.2},
  {1.2, 3.8, 2},
  {3.6, 3.4, 3.6},
  {3, 1.6, 3.2},
  {3, 0.6, 1.8},
  {5, 1, 2.6},
  {5.4, 3.8, 4.2},
  {6, 4.2, 5.4},
  {9.4, 7.4, 10.2},
  {5.8, 6.8, 8.2},
  {0.4, 1.6, 1},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1, 0.2, 0.2},
  {1, 0, 1.2},
  {0.6, 0, 0},
  {0.6, 0, 0},
  {0, 0, 0},
  {0, 0.4, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0.6, 0.2},
  {0.6, 0.8, 0.8},
  {0.2, 1, 0.4},
  {0.2, 0.4, 0.4},
  {0, 0, 0.2},
  {0, 4.2, 1},
  {0.2, 1.4, 1.2},
  {0, 3, 0.6},
  {0, 1.4, 0},
  {0, 1.8, 0},
  {0, 2, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.4, 0},
  {0.2, 0.2, 1.8},
  {1, 0.6, 1.4},
  {0.6, 0, 1.2},
  {1.8, 0, 0},
  {2.4, 0, 0},
  {2, 0, 1.8},
  {1.4, 0, 0},
  {6.8, 0, 1.6},
  {8, 0, 6.4},
  {4.2, 0, 3},
  {2, 0, 1.8},
  {5.6, 0, 1},
  {7, 0, 1.8},
  {1.4, 0, 1},
  {1.2, 0, 0.8},
  {0, 0, 0},
  {0, 0, 0},
  {0.8, 2.8, 1},
  {1.2, 2, 2},
  {3.6, 0.4, 3.2},
  {0.8, 0.4, 1.4},
  {1, 0.2, 0.4},
  {0.2, 0.4, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0.4},
  {0.2, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1.2, 0.4, 0},
  {0, 0.2, 0.4},
  {0.2, 0, 0},
  {0.4, 0.2, 0},
  {0, 0, 0.2},
  {0.6, 0, 0.6},
  {2.4, 0, 0.2},
  {3.8, 0, 4},
  {2.8, 0, 2},
  {0, 0, 0.8},
  {0, 0, 0.2},
  {0.2, 0, 0},
  {0.6, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0.2, 0.6},
  {1.6, 0.6, 0.8},
  {2.4, 2, 1.4},
  {0.4, 1.8, 0.8},
  {0, 1.2, 0.8},
  {0, 1.6, 0},
  {0, 2, 0},
  {0, 0.4, 0},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.6, 0, 0.4},
  {0, 0.2, 0.4},
  {0.2, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1, 0, 0},
  {1.4, 0.2, 0.4},
  {1.2, 1.4, 0.8},
  {0.4, 0.6, 0.6},
  {0.2, 0.2, 0.4},
  {0, 0, 0.4},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.6, 0.4, 0},
  {0, 0, 0.4},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0.4, 0, 0.6},
  {0.6, 0.2, 0.2},
  {0.2, 0, 0.2},
  {0.2, 0, 0},
  {0.2, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.4, 0, 0},
  {0.2, 0, 0.4},
  {0, 0.4, 0.4},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.6, 0, 0},
  {1, 0, 0},
  {0.8, 1.2, 1.8},
  {0.8, 1, 1.2},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0.4, 0, 0.4},
  {0.2, 0, 0.2},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.6, 0.4, 0.8},
  {0.2, 1, 0},
  {0.8, 0.6, 0.2},
  {1.2, 1.2, 0.6},
  {0.2, 0.4, 0},
  {0, 0, 0},
  {0.8, 0, 0},
  {0.6, 0.8, 0.8},
  {0.8, 0.8, 0.6},
  {1.2, 1.2, 1.8},
  {2.8, 2.6, 1.8},
  {3, 3.4, 4.2},
  {1.4, 3.2, 4.2},
  {0.2, 2.4, 1.6},
  {0, 1.2, 0.8},
  {0.2, 0.8, 0.6},
  {0.4, 0.2, 1},
  {0, 1.2, 0.6},
  {0, 0.4, 0.4},
  {0.2, 0, 0.4},
  {1.6, 0.4, 0.8},
  {2.2, 1, 1.4},
  {2.4, 2.2, 2.8},
  {1.2, 0.6, 2},
  {1.4, 0.4, 1.8},
  {1.6, 0.4, 3},
  {0.2, 0.2, 1.2},
  {0.2, 1, 0.4},
  {0.8, 0.8, 0},
  {0.2, 0, 0.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.8, 0, 0},
  {1.8, 0, 0.2},
  {0.4, 0, 0.6},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.6, 0, 0},
  {0.8, 0.2, 0.2},
  {0.6, 0.6, 0},
  {0.4, 0.8, 0.6},
  {0.4, 0.2, 0.2},
  {0.2, 0.4, 0.2},
  {0.2, 0.2, 0},
  {0.2, 0.6, 0.2},
  {0.2, 1.2, 0.4},
  {0, 0.8, 0.4},
  {0.2, 1, 0.2},
  {0, 1, 0.4},
  {0, 0.6, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0.8, 0.4, 0.6},
  {1, 1, 1},
  {1.8, 1, 1.6},
  {1.8, 0.6, 1.8},
  {1.4, 0.6, 1.8},
  {0.6, 0.4, 1.2},
  {0, 0, 0.2},
  {0.4, 0, 0.6},
  {0.2, 0.2, 0.8},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0.6, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1, 0, 0.8},
  {0.6, 0.4, 1.6},
  {2.2, 0.6, 2},
  {1.4, 1, 2.4},
  {1.6, 0.4, 2.2},
  {0.8, 0, 1.4},
  {0, 0.2, 1.4},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.8, 0.2, 0},
  {2, 1.8, 0.4},
  {1.4, 2.2, 1.2},
  {0.2, 1, 1},
  {0, 1, 0.4},
  {0.2, 1, 0.6},
  {0.6, 0.8, 1.2},
  {0.2, 0.6, 1},
  {1.6, 0.8, 2},
  {3.2, 1.2, 4.2},
  {3, 3.2, 4.6},
  {2.4, 3, 3.6},
  {5.2, 3.2, 4.4},
  {4, 4.8, 7.2},
  {5, 4.2, 5.6},
  {1.6, 2.6, 4.2},
  {0.6, 1.6, 1.6},
  {0.4, 1.4, 1.6},
  {4, 0.6, 3.2},
  {0.6, 3.8, 1.6},
  {0.2, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0.2, 0},
  {0.2, 0.2, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0.2, 1.4, 0.4},
  {0.2, 0.8, 0.4},
  {0.4, 0.2, 0.2},
  {1.4, 3, 2.6},
  {0.4, 2, 0.6},
  {0.4, 0.4, 0},
  {0, 0.2, 0.2},
  {0.4, 0.8, 1},
  {1.8, 3.2, 2.4},
  {0.4, 3, 0.6},
  {0.2, 0.2, 0},
  {0, 0.6, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.8, 0, 0},
  {0.8, 0, 0},
  {0.2, 0.2, 1.8},
  {0.2, 0.2, 0.4},
  {0, 0, 0.4},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.2, 0, 0},
  {0.4, 0, 0},
  {0.2, 0, 0.2},
  {0.2, 0, 0.2},
  {0.2, 0, 0},
  {0, 0, 0.4},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.4, 0, 0.2},
  {0, 0, 0.2},
  {0, 0.2, 0.6},
  {0, 0, 0.6},
  {0, 0, 0.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.6, 0, 0},
  {0.2, 0, 0.4},
  {0.2, 0, 0},
  {1, 0, 0},
  {0.8, 0, 0.6},
  {0.8, 0, 0.2},
  {1, 0, 0},
  {1.4, 0, 0},
  {2, 0, 0.2},
  {2, 0.2, 0},
  {2.8, 0, 0},
  {2.2, 0, 0},
  {2.2, 0.2, 0},
  {1.6, 0, 0},
  {0.2, 0, 0},
  {0.4, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0, 0.2, 0.2},
  {0.2, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0.2, 0},
  {0.6, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.6, 0, 0.8},
  {1.2, 0.6, 1.2},
  {0.8, 0.8, 1.6},
  {0.8, 0.6, 1.4},
  {0.4, 0.4, 1.2},
  {0.6, 0.2, 0.8},
  {1.6, 0, 1.2},
  {1.4, 0.2, 2},
  {0.6, 0.6, 1.8},
  {1, 0.6, 1.2},
  {1, 0.6, 2.4},
  {1.2, 0.4, 2},
  {1.4, 0.4, 2.6},
  {1, 0.4, 1.6},
  {0.6, 0.2, 1.8},
  {0.4, 0.6, 0.6},
  {0.6, 0.2, 1},
  {0.8, 0.2, 1.8},
  {0.8, 0.2, 1.8},
  {1.8, 0, 1.2},
  {2.4, 0.6, 2.4},
  {0.6, 0.8, 2},
  {0.8, 0.8, 2.4},
  {1, 1.6, 2.4},
  {0.4, 1, 1.4},
  {0.6, 0.2, 1.4},
  {0.4, 0.4, 1.6},
  {1.2, 0.6, 0.6},
  {0.2, 0.8, 1.4},
  {0.4, 0, 0.4},
  {0.6, 0.6, 1.2},
  {0, 1.4, 1},
  {1.2, 0.6, 0.8},
  {0.4, 0.6, 1.8},
  {0, 0.4, 1.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0.2, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.6, 0, 0},
  {0.2, 0.2, 0},
  {0.4, 0.2, 0.2},
  {1.6, 0.2, 0.4},
  {1, 1.8, 2},
  {1.6, 1.8, 2.6},
  {3, 4.8, 5},
  {4.4, 5.6, 7.6},
  {3.6, 2.6, 3.6},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0.2, 0},
  {0.2, 0.6, 0},
  {0.4, 0.4, 0.6},
  {0.2, 0.8, 2},
  {0, 0.6, 1.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0.2, 0, 1.2},
  {0, 0, 2.2},
  {0, 0, 0.2},
  {0.6, 0, 1},
  {1.6, 0.2, 2},
  {2.8, 1.8, 4},
  {3, 2, 3.4},
  {2.8, 2.8, 5.2},
  {1.6, 1.8, 2.8},
  {1, 2, 2},
  {0, 1.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0.2, 1.8},
  {0.2, 0.6, 0.6},
  {0, 1.2, 1.4},
  {0.2, 0, 1.6},
  {0.8, 1, 1.2},
  {1.8, 1.4, 0.2},
  {0.8, 0.4, 0.6},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0.2},
  {0.6, 0, 0.2},
  {0.2, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0.2},
  {0.2, 0.2, 0},
  {0.2, 0, 0.2},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0.6, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.6},
  {0, 0, 1.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1.4, 0, 0},
  {0.8, 0, 0},
  {0.4, 0, 0},
  {0.4, 0, 0},
  {1, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0.4},
  {0, 0, 0.6},
  {0, 0, 0.2},
  {0.2, 0, 0.2},
  {0.2, 0, 0.2},
  {0.2, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.6, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0.2, 0, 0.2},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 1.8, 1.4},
  {0, 0, 0.2},
  {0, 0, 1},
  {0, 0, 0.2},
  {0, 0, 0},
  {0.4, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1.8, 0, 0},
  {2.6, 0, 0.2},
  {3.4, 1.2, 1.4},
  {2.6, 2.2, 2.2},
  {3.4, 3.6, 3},
  {2.6, 3.6, 5},
  {3.2, 2.6, 4.4},
  {4.8, 4.6, 4.6},
  {3.2, 6, 3},
  {0, 5, 0},
  {0.2, 0.2, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.4, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {1.8, 0, 0.2},
  {1.6, 0.6, 1},
  {2, 2.2, 1.6},
  {0.8, 2.2, 1.4},
  {0, 0.4, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.8, 0, 0.4},
  {0.4, 0.2, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0.4, 0, 0},
  {0.4, 1.2, 0.4},
  {1, 0.6, 0.2},
  {0.6, 0.6, 0.2},
  {0.8, 1, 0.8},
  {1.6, 0.8, 1.6},
  {2.6, 0.8, 1.4},
  {2, 4.8, 2.2},
  {6.8, 0.6, 0.2},
  {7.2, 0, 0.6},
  {8.8, 7.4, 1.4},
  {11.2, 5.2, 9.8},
  {13.6, 0.6, 10.4},
  {2, 0, 2.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.6, 0},
  {0, 0.6, 0},
  {2.4, 0, 0.6},
  {0.6, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0.2, 0.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1.2, 0, 0},
  {1.8, 1.4, 0.6},
  {0.4, 2, 1},
  {1.4, 2.4, 1.8},
  {0.2, 0.4, 0.2},
  {1, 0.8, 0.4},
  {0.2, 0.4, 0.4},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.4, 0},
  {0, 1.2, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0.2, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0.2},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.4, 0.2, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.6, 0.4, 1.2},
  {0.2, 2.6, 2.6},
  {1, 0.8, 2.8},
  {0, 1.6, 5.4},
  {1.4, 1.6, 2.6},
  {1.2, 4.6, 3.4},
  {2.8, 5.8, 5.6},
  {6.2, 3.6, 4.4},
  {1.2, 4, 3.6},
  {3, 1.6, 1.4},
  {0, 0.4, 1},
  {0.6, 0.8, 0},
  {0.2, 0, 0},
  {0, 0.2, 0},
  {0, 0.6, 0},
  {0, 1.4, 0},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1.2, 1, 0.6},
  {0.6, 0.8, 1.2},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1.2, 0, 0},
  {0.4, 0, 0},
  {0.2, 0, 0.2},
  {0.6, 0, 0.2},
  {1, 0, 0},
  {0.6, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0.2, 0.8, 0.2},
  {0, 0.2, 1.2},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0.2, 0},
  {0.2, 0, 0},
  {0.2, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.2, 0, 0},
  {0, 0.6, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0.2},
  {0, 0.2, 0.2},
  {0.2, 0.2, 0.6},
  {0.2, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {2, 0, 0},
  {2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1.6, 0, 0},
  {5, 0, 0.4},
  {1, 0, 2},
  {0, 0, 0.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 1, 0.4},
  {1.6, 4, 3.4},
  {3.2, 9.4, 2},
  {3.6, 5.2, 3.8},
  {5.2, 3, 3.8},
  {1.8, 3.2, 2.2},
  {0, 1.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0.4},
  {0.6, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.6, 0},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0.2, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0.2, 0},
  {0, 0.8, 0},
  {2.6, 0, 0},
  {3.8, 2.2, 3.4},
  {1.2, 2.2, 3.6},
  {0.6, 2, 4.6},
  {5.6, _, 2.8},
  {4.2, 3.8, 6.2},
  {0.2, 1.2, 5.4},
  {0.2, 1.8, 1.8},
  {0.2, 2.2, 0},
  {3.4, 0.4, 0.4},
  {4, 3.6, 3.8},
  {2.4, 3.2, 2},
  {1.2, 0.6, 0.2},
  {0.2, 0.4, 0.4},
  {0.8, 0, 0.2},
  {2.8, 0.2, 1},
  {1.8, 0.4, 1.2},
  {1, 0.2, 1.4},
  {0.8, 0, 0.4},
  {1.6, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 4.2, 1},
  {0, 5.8, 0.8},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.6, 0, 0},
  {0, 0, 0},
  {1.8, 1, 0},
  {4, 2, 1},
  {5, 1.2, 2},
  {0.4, 0.4, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.6},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 1.8, 0.2},
  {0, 0.4, 1.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0, 0, 0.8},
  {0.2, 0, 0.2},
  {0.2, 0.6, 0},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 4},
  {0, 0, 1.8},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.8},
  {0.8, 2.2, 3.4},
  {0.2, 0.8, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 2.6, 0},
  {0, 1.4, 0.8},
  {0, 5.6, 1.4},
  {10.6, 0.2, 3},
  {0, 0, 0},
  {0.4, 2.8, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 2, 0},
  {0, 0, 0},
  {0.2, 0.2, 0},
  {1.8, 0, 0.4},
  {0.8, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {3.4, 0, 2.6},
  {4.6, 0, 2.2},
  {2.4, 1.4, 0.4},
  {2.8, 0.2, 1.4},
  {0.6, 0, 1.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {2.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {4.8, 0, 0},
  {0.2, 0, 0},
  {2.8, 0, 0},
  {8.2, 0, 0.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 1.4, 0},
  {0, 1.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 2.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 3.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {3.6, 0, 0},
  {0.2, 7, 0.6},
  {1, 0.2, 0.2},
  {0, 0.6, 0.8},
  {6.8, 1.4, 3.8},
  {4.8, 2.8, 2.4},
  {1, 2, 0.6},
  {3.8, 0.8, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 2, 4.8},
  {0, 0, 0},
  {0, 0.4, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {3.6, 0, 0.2},
  {3.6, 0.2, 0},
  {0.6, 0.4, 3},
  {0, 0.6, 4.4},
  {0, 4.2, 9.8},
  {6, 3.8, 2},
  {0.8, 2.2, 2},
  {0.8, 2.2, 3.8},
  {7.2, 4, 2.2},
  {3.4, 6.4, 5.2},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {1, _, 3},
  {0.2, _, 0.4},
  {0.4, _, 2.6},
  {1.8, _, 5.2},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, _, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.8},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.6, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1.6, 0.2, 1},
  {2, 3.6, 3.2},
  {1.8, 6, 0.6},
  {0.4, 1, 1},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.6, 0, 0},
  {0.2, 0.2, 0.8},
  {0, 0, 1},
  {0, 0.2, 0.2},
  {0.2, 0, 0},
  {1.2, 0.2, 0},
  {2.8, 1.6, 0.2},
  {1.2, 1.4, 1},
  {0, 0.2, 1.2},
  {1, 0.2, 0.6},
  {0.6, 0, 0.8},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 1, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.6, 0, 0},
  {0.4, 0, 0.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.4},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 1},
  {0, 0, 0},
  {0, 0, 0},
  {2.4, 0, 0},
  {2.6, 0, 0},
  {0.4, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 4},
  {0.4, 0, 0.8},
  {0.8, 0, 0.4},
  {0, 0, 0.6},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 1.2},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 3.8, 0},
  {0, 0.6, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0.6, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 17},
  {0, 0, 1.4},
  {0, 0.2, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 13.4, 0},
  {0, 2.2, 0},
  {9, 3.2, 0},
  {0.2, 0, 0.6},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 2.8},
  {0, 0, 3.2},
  {0.8, 0, 4.8},
  {0.2, 2.2, 6.2},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0.6, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.4},
  {0.2, 0, 1},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {9, 0, 8.2},
  {0.2, 0, 0.2},
  {0.2, 0, 0.2},
  {0, 0, 0},
  {0, 0.6, 0.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {3.2, 1.2, 0.8},
  {3, 1.8, 2.8},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1.6, 0, 0.8},
  {6.2, 4, 1},
  {1.6, 1.8, 0.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 2.4, 0},
  {0, 0.2, 1},
  {0, 0.2, 0.2},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.6, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {1, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.6, 0},
  {0, 0.6, 0},
  {2.4, 0.2, 0},
  {5.2, 2.2, 2.2},
  {5, 2.6, 5.2},
  {3.8, 1.6, 3},
  {2.2, 1.4, 2.2},
  {3.8, 5.4, 3.2},
  {0.8, 2.2, 4},
  {2, 3.6, 3.8},
  {4.2, 7.6, 1.8},
  {10.6, 6.4, 6.8},
  {6.2, 8.8, 3.2},
  {5.8, 4, 9},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {1, 0, 0},
  {2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 1},
  {0, 0, 1.8},
  {0, 0, 0.4},
  {0, 0, 1},
  {0, 0, 1},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {3, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 3.8, 0},
  {0, 2.2, 0},
  {0.6, 0.2, 0},
  {0.4, 0, 0},
  {2, 0, 0},
  {0.2, 0, 0},
  {0.6, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 1.8, 0},
  {8.6, 0.6, 1.2},
  {3.2, 2.8, 0},
  {0, 2.2, 0.8},
  {1.6, 2.6, 1.6},
  {0.6, 0, 1.6},
  {1.4, 0, 0},
  {0, 0.2, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0.2},
  {0, 0, 10.6},
  {0, 0, 1},
  {0, 0.2, 0},
  {0, 8.4, 0},
  {2.8, 0, 0},
  {1.6, 0, 0},
  {0.2, 4.2, 0.2},
  {1, 5.2, 1.2},
  {3.4, 0.4, 2.2},
  {2.4, 0.2, 0},
  {0.2, 0.8, 0.2},
  {0.4, 0.4, 0},
  {0.4, 0.4, 0.8},
  {0.4, 0.6, 0.4},
  {0, 0.2, 0.6},
  {0, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1.8, 0, 2},
  {0, 2, 0.8},
  {2, 0, 1},
  {2.4, 0, 0.2},
  {0.8, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.8, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {3, 0, 0},
  {4.2, 1.8, 0.2},
  {0, 1.8, 0.8},
  {0, 0, 1.6},
  {0, 0, 0.2},
  {0, 0, 0.2},
  {0, 0, 0},
  {0.2, 0.6, 0.2},
  {0, 0.6, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.6, 0.2},
  {0, 2.2, 0},
  {0, 0, 0},
  {0.8, 0, 0},
  {0.6, 0.6, 0},
  {0, 0, 0},
  {0, 0, 0.4},
  {0, 0, 1.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {1, 0.6, 0},
  {0.4, 0.4, 1.2},
  {1.4, 3.2, 0.4},
  {1.6, 0.8, 2.6},
  {1.2, 4.4, 1.8},
  {0.4, 0.2, 3},
  {5.8, 2.2, 0},
  {11.6, 9.4, 3.2},
  {0.8, 7, 2.6},
  {2.4, 0.8, 0.6},
  {0.6, 0.2, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {1.8, 0.8, 0},
  {0.4, 1.2, 0},
  {3.4, 2.2, 0},
  {0.4, 4.4, 0},
  {0, 0, 0.6},
  {0.2, 0, 0},
  {0.4, 0, 0},
  {0, 0.2, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 1, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.6, 0, 0},
  {1.2, 0.2, 0},
  {0, 0, 0},
  {0, 0.4, 0},
  {0, 0.4, 0.4},
  {0.2, 0, 0.6},
  {3.6, 0, 0.6},
  {0.4, 0.6, 1.8},
  {2.2, 7.2, 2.2},
  {2.8, 4.6, 1},
  {0.4, 0.4, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0.8, 0, 0},
  {0.2, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {3.8, 0, 0},
  {0, 3.2, 0.2},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 1.2},
  {1.4, 4.2, 1.8},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 5.4, 0},
  {0, 1.6, 0},
  {0, 0, 0},
  {1, 0, 0},
  {0.2, 2, 0},
  {0.2, 0, 0},
  {0, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {1.6, 0, 0},
  {0, 0.2, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0.4},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.8, 0, 0.2},
  {0, 0, 0},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 5.4},
  {6.2, 13.8, 7},
  {2, 4, 7.2},
  {1.8, 2.6, 3.4},
  {0, 1.6, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 6},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0.6, 0.8, 0},
  {1, 0.6, 0.2},
  {0.2, 1, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0.6},
  {1.6, 0, 0.4},
  {0, 0, 0},
  {0.4, 0, 0},
  {0.2, 0, 0},
  {1.4, 0, 0},
  {0.6, 1.2, 0},
  {0.4, 1, 0.2},
  {1.2, 1.6, 0},
  {2.8, 3.4, 0.2},
  {3, 4.4, 1},
  {3.2, 5.4, 2.4},
  {5.8, 10.4, 3.6},
  {7.6, 15, 5},
  {6, 10.2, 9.8},
  {4, 12.2, 8.8},
  {4.4, 4.6, 7},
  {5.2, 8.2, 3.8},
  {0, 7.8, 4.2},
  {0, 1.4, 9.4},
  {0.4, 0.2, 1.6},
  {0.2, 0, 3},
  {0, 0.6, 3.4},
  {0, 2.6, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 1},
  {0, 0, 3},
  {0, 4.2, 1.6},
  {0, 3.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0.6},
  {0, 0.2, 0.8},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.8},
  {1.6, 1.8, 0.4},
  {1.2, 0, 0.4},
  {1.8, 1.4, 0.4},
  {3.6, 4, 1},
  {3.4, 1.4, 2.2},
  {0.2, 0.2, 0.6},
  {1, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {1, 1.2, 0},
  {0.4, 0.6, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.4, 0},
  {0.2, 0, 0},
  {0.2, 0.2, 0},
  {0, 0, 0},
  {0, 2, 0},
  {0, 0.4, 0},
  {0.2, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 1.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {1.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {_, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 1.2, 0.4},
  {0.8, 0, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 1.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.8, 0, 0},
  {2.8, 0.8, 0.6},
  {9.4, 4.2, 0.2},
  {2.6, 11.4, 1},
  {0, 1.4, 4.2},
  {0, 0, 1.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.2, 0.6, 0},
  {0.2, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.4},
  {0, 0, 1.6},
  {0, 0, 1.4},
  {0, 0, 1.4},
  {0, 0, 1.2},
  {0, 0, 0.4},
  {0, 0, 0.6},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0.2, 0},
  {1, 0.8, 0.2},
  {1.4, 0.4, 0},
  {1.6, 1.6, 0.2},
  {2.2, 1, 0.2},
  {0.4, 0.6, 0.2},
  {0, 0, 0.2},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.6, 0, 0},
  {1.6, 0, 0.2},
  {0.8, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.6, 0, 0},
  {1.8, 0.2, 0},
  {0.6, 0.6, 0},
  {0.4, 0.6, 0},
  {1, 0.4, 0},
  {1, 0.8, 0},
  {1.4, 1, 0},
  {1.4, 1, 0},
  {1, 2, 0},
  {2, 2.2, 0},
  {2.2, 4.6, 0},
  {0.4, 3.6, 0},
  {0.2, 2.8, 0},
  {0, 0.6, 0.2},
  {0, 0.2, 0},
  {0, 1, 0},
  {0.2, 0.8, 0.6},
  {1.2, 1, 1},
  {0.4, 2, 0.8},
  {1.2, 0.2, 0.6},
  {0.4, 0.8, 0.2},
  {0.6, 2.4, 0.4},
  {0, 0.6, 0.4},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.6, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, _},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, _},
  {0, 0, _},
  {0, 0, _},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.2},
  {0, 0, 0},
  {0.8, 0, 0},
  {5.4, 1.2, 0.2},
  {3.6, 2.6, 0.6},
  {0.4, 3, 1.8},
  {0, 0.4, 0.2},
  {0, 0.6, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 1.4, 0.6},
  {0, 0.6, 2.6},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0.4},
  {2.4, 0, 0.6},
  {0.2, 0.6, 0.6},
  {0, 0.4, 0.8},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0.4, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {2.6, 1.6, 2},
  {0, 0.6, 0},
  {0, 0, 0},
  {0, 0.6, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0, 0.2},
  {0.6, 0.4, 1},
  {0.6, 1, 0.6},
  {0.8, 1.4, 1.4},
  {1, 2.8, 0.8},
  {0.2, 1.4, 0.8},
  {0.4, 0, 0},
  {0, 0.4, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.4, 0, 0},
  {0.4, 0, 0},
  {1, 0, 0},
  {0.4, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {2, 0.4, 0.6},
  {0.2, 1.2, 0.8},
  {0.2, 2.4, 0.2},
  {0, 1.2, 0.8},
  {0, 0, 0},
  {0.6, 0.2, 0},
  {0, 0.6, 0.6},
  {0, 1, 0},
  {0, 2.2, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0.4, 0.4},
  {0, 0, 0.8},
  {0.4, 0.2, 2},
  {0, 0.2, 4.8},
  {0.8, 3.6, 4.6},
  {0, 2.2, 2.8},
  {0.6, 0.8, 0.4},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {1.4, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0.2},
  {0.2, 0, 0},
  {0.2, 1, 0.6},
  {0.2, 0.2, 0.2},
  {0, 0, 0},
  {0, 0.6, 0.2},
  {0.2, 2.6, 0.4},
  {0, 0.8, 1},
  {0, 0, 0.6},
  {0.2, 1.2, 1.2},
  {0, 0.8, 0.6},
  {0, 0, 0},
  {0, 0.4, 0.4},
  {0, 0, 0},
  {0, 0, 0.4},
  {0.2, 0, 0},
  {0, 0, 0.4},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 2},
  {0, 1.2, 0},
  {0, 0, 0},
  {0, 0, 0.4},
  {0.8, 0.4, 1},
  {0.4, 2.8, 2.4},
  {2.6, 4.2, 1.8},
  {3.8, 4.6, 4.6},
  {5, 5.2, 4.6},
  {6.8, 5.2, 5.4},
  {2, 4.8, 6.4},
  {2, 1.6, 1.4},
  {1.8, 0.2, 0.4},
  {1, 0.8, 0.6},
  {6, 2.2, 3.8},
  {1.2, 5.4, 5},
  {1.6, 0.6, 0.6},
  {0, 1.2, 1.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {3.6, 0, 0},
  {0.8, 0, 0},
  {0, 1.2, 0},
  {0, 4.4, 0},
  {0.8, 0, 0},
  {0.6, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.6, 0, 0},
  {1.6, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0.2, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.6, 0, 0},
  {0.8, 0.6, 0},
  {0.4, 0, 0},
  {0, 0, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.8, 0, 0},
  {1, 0, 0},
  {0.2, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.6, 0, 0},
  {0.4, 0, 0},
  {0.8, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 1.6, 0},
  {0.4, 3.4, 0.2},
  {0, 0, 1},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0.2, 0.2},
  {0, 0, 0.4},
  {0, 0, 0.2},
  {0, 1.8, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {1, 0, 0},
  {0.6, 1.2, 0.4},
  {1.2, 1.6, 0.6},
  {1.2, 3, 1},
  {0.2, 2.6, 2.8},
  {0, 0.8, 0.8},
  {1.2, 1.4, 0.2},
  {1.2, 2, 0.8},
  {2, 0.6, 2.8},
  {2, 3.8, 4.4},
  {3.2, 2.2, 2.6},
  {5.6, 3.4, 3.8},
  {3, 3.6, 4},
  {3.4, 2.4, 2.2},
  {1, 3.2, 1.8},
  {0, 0, 0.6},
  {1.4, 1.6, 0},
  {3.4, 3, 2.2},
  {6, 3, 3.6},
  {2.2, 1.4, 5.6},
  {2.6, 0.8, 3.6},
  {0.2, 2.8, 2},
  {0, 1.4, 6.2},
  {0.8, 0.6, 0.4},
  {2.4, 3.8, 1.6},
  {0, 2.8, 3},
  {0, 0.6, 0.4},
  {0, 0.2, 0.6},
  {0, 2.2, 1.6},
  {0, 1, 0.2},
  {0.8, 0, 0.2},
  {0, 2.2, 0},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0.4, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0.6, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.4, 0.4, 0},
  {1.2, 2.2, 1.2},
  {1.4, 3, 1},
  {2, 1.8, 1.2},
  {2, 1, 0.8},
  {0.8, 1.8, 0.4},
  {0, 0, 0.2},
  {0, 0, 0.2},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {1.8, 1.8, 0.4},
  {3, 3, 2.2},
  {2, 1.8, 3},
  {1.2, 1, 1.6},
  {1.6, 5.2, 1.2},
  {1.4, 5, 2},
  {0, 0.8, 0.6},
  {0, 0.2, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0.8, 0, 0},
  {1.4, 0.6, 0.8},
  {0.4, 1, 1},
  {0.2, 0.4, 0.8},
  {0.4, 1, 1.4},
  {0.8, 1.4, 0.8},
  {3, 3.2, 3},
  {0.4, 3.2, 2.4},
  {0.2, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0},
  {0, 0, 0} ;

 Temp =
  {-11, -9.9, -8.8},
  {-10.7, -10.5, -9.7},
  {-10.2, -10.9, -10.5},
  {-10.6, -11.3, -11.2},
  {-11.6, -11.5, -11.7},
  {-11.5, -12, -12.1},
  {-11.8, -12.5, -12.3},
  {-11.8, -12.9, -12.8},
  {-12.5, -12.8, -12.9},
  {-11.8, -12.2, -12.5},
  {-9.5, -10.3, -9.5},
  {-8.4, -7.8, -6.4},
  {-7.2, -6.2, -4.2},
  {-6.2, -5.2, -2.3},
  {-5.2, -3.8, -0.6},
  {-4.7, -2.6, 0.2},
  {-4.7, -1.7, -0.2},
  {-5, -2, -0.9},
  {-6.8, -3.5, -2.5},
  {-8, -4.9, -3.1},
  {-9.3, -5.9, -4.5},
  {-10, -6.7, -6.1},
  {-10.6, -7.5, -7.4},
  {-10.5, -8.3, -8.2},
  {-10.7, -8.8, -9.1},
  {-10.9, -9.4, -9.8},
  {-11.1, -9.5, -10.3},
  {-11.2, -9.6, -10.9},
  {-11.3, -9.5, -11.4},
  {-11.2, -9.6, -11.7},
  {-11.9, -10.1, -12.1},
  {-11.7, -10.6, -12.4},
  {-11.7, -10.4, -12.5},
  {-8.8, -9.1, -12.2},
  {-5.9, -7.7, -9},
  {-4.7, -4.7, -5},
  {-2.8, -3.7, -1.5},
  {-1.8, -1.7, 0.8},
  {-0.6, 0.3, 2.9},
  {-0.1, 1.6, 2.9},
  {-0.3, _, 2.3},
  {-1.3, _, 1.2},
  {-2.7, _, 0.3},
  {-4.7, _, -0.5},
  {-5, -2.8, -2.6},
  {-6.3, -3.2, -3.6},
  {-7.8, -3.7, -4.8},
  {-7.9, -4.8, -5.4},
  {-8, -5.4, -6.1},
  {-8.2, -6, -7},
  {-8.5, -6.3, -7.1},
  {-8.8, -6.4, -7.7},
  {-8.8, -6.8, -8.1},
  {-9.4, -7, -8.2},
  {-8.8, -7.4, -9.1},
  {-7.2, -7.4, -9.1},
  {-6.3, -6.9, -8.3},
  {-6.1, -6.1, -6.9},
  {-5.9, -5.4, -5.3},
  {-6.3, -4.8, -4.4},
  {-6.7, -5.1, -3.9},
  {-5.9, -6.1, -3.9},
  {-6.2, -5.7, -3.6},
  {-5.6, -5.5, -3.4},
  {-4.9, -5.2, -2.8},
  {-4.9, -5, -2.8},
  {-4.7, -5.2, -3.2},
  {-5.3, -5.4, -3.5},
  {-5.4, -5.5, -3.5},
  {-5.5, -5.1, -3.6},
  {-5.7, -5, -3.7},
  {-5.4, -5.1, -3.7},
  {-5.4, -5.2, -3.7},
  {-6.7, -5.1, -4.4},
  {-7.8, -5.2, -8.5},
  {-8.4, -5.1, -7.6},
  {-8.4, -5.2, -6.2},
  {-8.7, -6.1, -5.9},
  {-8.8, -6.7, -5.9},
  {-8.7, -6.5, -5.5},
  {-8, -6.1, -5.6},
  {-6.4, -5.1, -5.6},
  {-2.8, -5.8, -5.5},
  {-2, -3, -4.7},
  {-0.8, -1.6, -2.9},
  {0.1, 0.5, 0.5},
  {1.9, 2.9, 1.9},
  {1.9, 3.7, 4.7},
  {2.5, 4.4, 6.7},
  {1.8, 4.1, 3.7},
  {-0.7, 0.8, 2.5},
  {-2.6, -0.2, -0.2},
  {-2, -0.5, -1.2},
  {-2.2, -0.5, -1.5},
  {-2.5, -0.7, -2.2},
  {-2.8, -1, -2.2},
  {-2.6, -1.5, -3.2},
  {-2.4, -2.4, -4.1},
  {-3.6, -2.6, -5.5},
  {-4.9, -2.9, -5.9},
  {-5.1, -3.3, -6.4},
  {-4.2, -4, -6.8},
  {-5.4, -4.4, -7.3},
  {-6.3, -5, -8.9},
  {-6.7, -4.8, -9.7},
  {-4.8, -4.3, -7.9},
  {-1.9, -3.4, -5.1},
  {-0.9, -1.2, -2.3},
  {-0.7, 0.8, 0.7},
  {0.3, 2.3, 4.5},
  {0.8, 2.8, 5.3},
  {0.3, 3.4, 4.2},
  {-1.2, 3.3, 3.2},
  {-1.1, 2.1, 2.6},
  {-2.1, 0.6, 2.3},
  {-2.5, -0.1, 1.2},
  {-3, -0.3, -0.8},
  {-3.3, -0.9, -2.9},
  {-4.2, -1.6, -3.9},
  {-5, -1.9, -4.7},
  {-5.3, -2.5, -5},
  {-5.3, -3.2, -6.6},
  {-5.8, -3.9, -7.4},
  {-6.1, -4.2, -8.2},
  {-6, -4.5, -8.2},
  {-6, -5, -8.6},
  {-6.5, -5.5, -9.6},
  {-6.9, -5.5, -10},
  {-6.6, -5.3, -10.4},
  {-4.4, -4.6, -9.4},
  {-1.4, -3.3, -6.6},
  {-0.6, 0.4, -3},
  {0.5, 1.8, 0.9},
  {1.3, 2.9, 3.8},
  {2.1, 3.6, 5.4},
  {1.7, 3.8, 5.4},
  {1.6, 3.5, 5},
  {0.3, 2.3, 3.7},
  {-0.6, 1.1, 3.1},
  {-1, -0.1, 3.6},
  {-1.7, -1.2, 3.3},
  {-2, -1.7, 2.5},
  {-3.3, -2.3, 1.7},
  {-4.5, -3, 0.7},
  {-5.4, -3.7, -2.4},
  {-5.7, -4.2, -3.5},
  {-6.2, -4.9, -4.1},
  {-6.6, -5.1, -5.6},
  {-6.8, -4.9, -7.3},
  {-7.8, -5, -8.3},
  {-9, -5.3, -8.8},
  {-8.8, -6.2, -10.1},
  {-8.4, -6.1, -10.1},
  {-6.8, -5.2, -9.4},
  {-4.1, -3.5, -6},
  {-3, -2.1, -2.4},
  {-2, -0.9, 0.8},
  {-0.5, 0.3, 1.9},
  {0.2, 1.4, 3},
  {0.9, 2, 3.6},
  {1.1, 2, 4.1},
  {0.6, 1.4, 4.5},
  {-0.8, 0.5, 4},
  {-2, -0.2, 2.9},
  {-2.5, -0.8, 1.7},
  {-3.2, -1.1, 2.2},
  {-4.1, -1.4, 0.6},
  {-4.8, -1.9, -2.1},
  {-5.5, -2.4, -3.8},
  {-6.1, -2.4, -5.3},
  {-5.4, -2.8, -5.8},
  {-4.5, -3.4, -5.8},
  {-4.4, -4, -6.7},
  {-5, -4.6, -7.9},
  {-5.5, -4.6, -8.2},
  {-6.7, -5, -8.9},
  {-6.4, -5.2, -9.2},
  {-3.7, -4.3, -8.4},
  {-0.5, -2.8, -5.1},
  {0.8, -0.1, -1.8},
  {2, 3.3, 1.4},
  {3.2, 5.1, 4.4},
  {4, 6.4, 6.8},
  {4.6, 7.1, 8.3},
  {4.6, 7.5, 8.9},
  {4.4, 7.7, 7.6},
  {2, 6.1, 5.9},
  {-0.2, 3.6, 2.4},
  {-0.6, 2.4, 0.2},
  {-0.6, 2, -1},
  {0, 1.5, -2},
  {0, 1, -2.5},
  {-0.4, 0.4, -3.2},
  {0, 0.3, -3.9},
  {-0.7, 0.3, -4.4},
  {-0.7, 0.2, -4.7},
  {-1.4, 0, -5.1},
  {-2.1, 0.3, -5.4},
  {-2.3, 0.8, -6},
  {-1.9, -0.1, -6},
  {-0.9, 0, -5.6},
  {0.7, 1.2, -4.2},
  {2.5, 2.7, -1.7},
  {3.6, 5.1, 1.4},
  {4.8, 6.5, 4.7},
  {6, 7.8, 8.7},
  {7, 8.8, 10.5},
  {7.3, 9.1, 11.8},
  {7.4, 9, 11.4},
  {6.4, 8.7, 9.9},
  {4.3, 6.4, 8.1},
  {2.2, 5.5, 5},
  {1.3, 4, 2.8},
  {2.2, 3.1, 2.9},
  {1, 2.7, 1.7},
  {0.1, 2.3, -0.1},
  {-1.2, 2.1, -0.9},
  {-0.6, 1.6, -2},
  {-1.3, 0.9, -2.5},
  {-2.1, 0.4, -3.1},
  {-1.7, 0.1, -3.6},
  {-1.6, -0.1, -4.2},
  {-2.6, -0.7, -4.6},
  {-2.4, -0.9, -5.1},
  {-2.4, -0.4, -5.2},
  {0, 1, -4.5},
  {2.8, 3, -1.3},
  {3.9, 5, 2.2},
  {5.1, 6.8, 6.1},
  {6.4, 7.8, 9.4},
  {6.8, 8.8, 10.3},
  {7.3, 9.4, 11.4},
  {7.9, 9.5, 12.4},
  {7.5, 9, 10.9},
  {4.2, 7.6, 7.6},
  {3.9, 5.2, 3.5},
  {2.4, 4, 1.9},
  {1.2, 2.8, 0.8},
  {-0.4, 1.3, -0.4},
  {-0.8, 0.6, -1},
  {-2.1, -0.4, -1.6},
  {-2.3, -1, -2.1},
  {-3, -1.4, -2.6},
  {-3.1, -1.7, -3},
  {-2.9, -2.2, -3.5},
  {-2.6, -2.6, -3.6},
  {-2.5, -2.9, -4},
  {-2.3, -3.2, -4.1},
  {-2.2, -2.2, -3.4},
  {-2.1, -1.9, -2.4},
  {-2, -0.1, -1.3},
  {-1.5, 1.8, 0.1},
  {0.1, 2.8, 3.3},
  {1.6, 4.2, 4.6},
  {3.6, 5.4, 5.9},
  {4.9, 6.3, 7.4},
  {5, 5.9, 8.3},
  {4.9, 5.6, 8.6},
  {4.4, 5.8, 8.3},
  {3.7, 4.7, 6.7},
  {3.2, 4, 3.9},
  {2.5, 3.5, 2.8},
  {2, 2.9, 1.6},
  {2, 2, 1},
  {2.1, 1.4, 0.3},
  {2.1, 0.8, -0.2},
  {2.5, 1.7, -0.9},
  {2.8, 1.9, -1.5},
  {2.8, 1.1, -1.9},
  {2.6, 0.4, -2.2},
  {2.5, 0.1, -2.4},
  {2.2, -0.1, -2.9},
  {2.3, -0.1, -2.8},
  {3, 0.3, -2.1},
  {4.4, 2.3, 0.3},
  {5.3, 4.2, 3},
  {6.2, 6.6, 5.3},
  {7, 8.5, 9.9},
  {7.4, 9.8, 10.6},
  {7.6, 10.2, 10.6},
  {7.2, 10.2, 10.4},
  {6.9, 9.5, 10.1},
  {5.9, 8.1, 9.4},
  {5.1, 6.9, 8.6},
  {4.5, 6.3, 6.7},
  {4, 5.6, 4.3},
  {3.5, 4.4, 3.2},
  {2.6, 3.1, 1.9},
  {0.8, 2.5, 1},
  {0.5, 3.2, 0.1},
  {0.9, 3, -0.4},
  {0, 2.9, -0.1},
  {-0.1, 2.3, -0.7},
  {0.2, 1.8, -1.5},
  {-0.1, 1.3, -2.2},
  {-0.9, 1.2, -2.6},
  {-0.3, 1, -2.8},
  {1.7, 1.4, -2.2},
  {4, 3, 1.9},
  {5.2, 4.8, 6.4},
  {5.8, 6.2, 8.9},
  {6.8, 7.4, 9.7},
  {7.6, 8.8, 10.9},
  {7.6, 9.7, 11.8},
  {7.3, 10.2, 10.5},
  {6.7, 10, 10},
  {5.7, 7.9, 8.8},
  {3.8, 6, 6.7},
  {2.8, 5.3, 4.2},
  {1.6, 4.7, 2},
  {1.3, 3.9, 1.4},
  {1.4, 3.4, 0.5},
  {1.7, 2, -0.2},
  {-0.3, 1.4, -0.9},
  {-0.6, 0.6, -1.2},
  {-0.3, 0.1, -1.6},
  {-0.3, 0.2, -1.5},
  {-0.5, 0.4, -1.5},
  {-1.1, 0.2, -1.8},
  {-1.1, 0.2, -2.1},
  {0.7, 0.6, -2},
  {2.6, 1.6, -0.5},
  {4.1, 3.3, 1.6},
  {4.8, 4.6, 4.5},
  {5.9, 6.6, 7.9},
  {7, 8.4, 10.3},
  {7.5, 9.6, 11},
  {7.8, 10.2, 10.2},
  {7.2, 9.9, 9.4},
  {6.7, 8.9, 9.3},
  {5, 7.5, 8.6},
  {4.1, 6.2, 6.2},
  {2.2, 5, 4},
  {1.4, 5, 2.3},
  {1.1, 4.3, 1.3},
  {0.8, 3.7, 0.7},
  {1.1, 3.3, 0.3},
  {2.2, 3.1, 0.3},
  {2.4, 3, 0.2},
  {2, 2.9, -0.1},
  {1.3, 2.5, -0.2},
  {0.6, 2.2, -0.6},
  {0.9, 1.8, -1.2},
  {0.9, 1.6, -1.4},
  {1, 1.6, -1.5},
  {3.2, 3, -0.3},
  {5.9, 5.2, 2.7},
  {6.9, 7.3, 6},
  {8.2, 8.1, 9.6},
  {9.4, 10.1, 12.5},
  {10.5, 12.1, 14.4},
  {10.7, 13.5, 14},
  {10.9, 13.4, 13},
  {9.7, 12.5, 12.7},
  {7.6, 10.7, 11.4},
  {5, 9, 8.9},
  {3.9, 7.7, 6},
  {3.7, 7.4, 4.2},
  {3.1, 5.8, 2.8},
  {2.9, 5.3, 1.7},
  {2.7, 4.8, 1.4},
  {2.5, 4.3, 0.4},
  {2.2, 3.9, 0.4},
  {2.6, 3.9, -0.2},
  {2.6, 3.7, -0.3},
  {1.9, 3.6, -0.8},
  {1.6, 3.6, -1},
  {2.5, 2.7, -1.1},
  {2.8, 3, -1.1},
  {5.8, 3.9, -0.3},
  {9, 7.4, 2.8},
  {9.9, 8.8, 6.7},
  {10.7, 10, 11.4},
  {12.1, 12.6, 14.8},
  {13.5, 14.4, 16.6},
  {13.7, 15.9, 17.3},
  {13.4, 16.7, 16.9},
  {13.1, 15.4, 15.8},
  {11.5, 13.2, 14.1},
  {8.2, 11.1, 10.2},
  {6.7, 10.6, 7.2},
  {6.2, 9.2, 5.1},
  {5.2, 7.8, 3.7},
  {4.9, 7, 2.6},
  {4.7, 6.4, 1.7},
  {3.9, 5.8, 1.2},
  {4, 5.7, 0.9},
  {4, 5.5, 0.2},
  {3.2, 4.9, 0.1},
  {3.5, 4.7, -0.2},
  {3.7, 4.6, -0.5},
  {3.8, 4.3, -0.9},
  {4.1, 4.3, -0.6},
  {7.3, 5.7, 0.4},
  {10.1, 8.3, 4.1},
  {11.3, 10.7, 8.1},
  {13.5, 11.7, 12.5},
  {14.6, 13.9, 16.2},
  {15.2, 15.9, 18.8},
  {16.1, 17.2, 19.2},
  {15.2, 17.9, 18.7},
  {15, 16.9, 18.2},
  {12.8, 15.7, 15.8},
  {9.6, 12.7, 12.1},
  {9.1, 11.6, 8.5},
  {8.1, 10.5, 6.5},
  {7.4, 9.6, 5.1},
  {7, 9, 4.1},
  {6.9, 8.3, 3.4},
  {6.8, 8.2, 2.7},
  {6.1, 8.2, 1.9},
  {6.5, 7.3, 1.5},
  {6.4, 7.3, 0.8},
  {6.1, 7.1, 0.7},
  {6.5, 6.7, 0.2},
  {6.1, 6.5, 0.1},
  {7.2, 8.2, 0},
  {12, 10.5, 1.4},
  {14, 12.7, 5.5},
  {15.3, 15.2, 11.1},
  {16.5, 17.5, 16.4},
  {18, 19, 20.7},
  {18.9, 20.3, 23.1},
  {19.1, 21.1, 23.9},
  {18.6, 21.5, 22.2},
  {17.2, 21.7, 20.7},
  {15.5, 19.7, 17.2},
  {13, 15.6, 13.7},
  {11.3, 13.5, 10.1},
  {10, 12, 8},
  {9.8, 11.5, 6.6},
  {10.3, 10.9, 5.2},
  {9.4, 10.6, 4.3},
  {9.1, 10.8, 3.4},
  {8.4, 10.3, 2.6},
  {8.4, 10, 2.3},
  {8.2, 9, 2},
  {8.7, 9, 1.5},
  {8.4, 8.8, 1.1},
  {8.9, 7.7, 1.1},
  {8.9, 7.2, 1.1},
  {13, 9.5, 3},
  {15.2, 14.4, 7.5},
  {16.2, 17.2, 13},
  {17.8, 18.4, 18.4},
  {19.2, 19.8, 21.7},
  {19.7, 20.7, 23.6},
  {20, 21.4, 24.6},
  {19.8, 21.5, 23.5},
  {19.1, 21.5, 20.3},
  {16.1, 20.1, 18.4},
  {13.5, 17.5, 14.8},
  {12.6, 16.1, 12},
  {12.4, 15.3, 10.3},
  {11.8, 14.3, 8.2},
  {10.3, 13.6, 6.7},
  {10.9, 13.1, 5.8},
  {9.4, 12.1, 4.7},
  {8.5, 11.4, 4.2},
  {7.9, 10.8, 3.4},
  {7.4, 9.8, 3},
  {6.2, 8.7, 2},
  {6.1, 8.1, 2.1},
  {6.2, 7.3, 1.4},
  {7.1, 7.6, 1.5},
  {8.2, 8.7, 3.6},
  {10, 10.5, 7.1},
  {10.1, 12, 12},
  {10.9, 13.3, 13.8},
  {11.8, 13.8, 14.6},
  {11.4, 13.6, 14.1},
  {10.2, 13.7, 13.6},
  {10.3, 13.3, 13.3},
  {9.2, 12.5, 13},
  {7.8, 10.7, 12},
  {6.7, 8.9, 10.8},
  {6.3, 7.9, 8.9},
  {5, 7.1, 6.4},
  {3.7, 6.9, 5.2},
  {3.8, 6.7, 4.9},
  {4.7, 6.7, 5.2},
  {5.2, 6.8, 5.3},
  {5.4, 6.9, 5.7},
  {5.4, 6.8, 5.6},
  {5.5, 6.7, 5.6},
  {5.4, 6.5, 5.5},
  {5.1, 6.3, 5.5},
  {4.9, 6, 5.5},
  {5.5, 6.1, 5.8},
  {5.6, 6.7, 6.2},
  {6.2, 7.2, 7.2},
  {6.7, 7.7, 8.4},
  {7.3, 8.8, 9.7},
  {8.4, 10.8, 11.3},
  {9.8, 12.4, 13.7},
  {10.5, 13.2, 15},
  {10.2, 13.3, 13.3},
  {8.4, 11.8, 12.5},
  {7.1, 10, 11.3},
  {6.2, 8.2, 9.6},
  {4.7, 6.6, 7.7},
  {3.6, 6.5, 5.9},
  {3.1, 6.5, 4.3},
  {2.9, 5.7, 3.2},
  {2.6, 4.9, 2.4},
  {2.4, 4.6, 1.8},
  {2.1, 4.2, 1.2},
  {2.2, 3.9, 0.8},
  {2.2, 3.5, 0.5},
  {1.8, 3.2, 0},
  {2, 2.9, -0.4},
  {4.1, 2.7, -0.2},
  {5.4, 3.7, 0.7},
  {5.9, 5.5, 2.5},
  {6, 6.5, 4.2},
  {6.2, 7.8, 6},
  {6.1, 9.1, 7.6},
  {6.7, 9.8, 8.8},
  {7.7, 10.8, 10.4},
  {8.1, 10.8, 11.7},
  {8.5, 10.8, 13.1},
  {7.6, 10.5, 12.5},
  {6.6, 8.9, 11.1},
  {6.1, 7.7, 10},
  {6.2, 7.7, 8.6},
  {6.1, 7.4, 7.2},
  {5.8, 7.3, 6.5},
  {5.5, 6.4, 5.8},
  {5.6, 6.3, 5.6},
  {5, 6, 4.9},
  {4.6, 5.5, 3.8},
  {4.1, 5.3, 3.4},
  {3.6, 5.1, 2.9},
  {3.2, 4.8, 2.4},
  {3.2, 4.6, 2.2},
  {4.1, 4.8, 2.3},
  {5.3, 5.9, 3.1},
  {6.3, 7, 5},
  {7.9, 8, 8.2},
  {8.4, 9.2, 10.9},
  {8.5, 11, 12.2},
  {8.4, 12.3, 12.2},
  {8.7, 12.3, 12.1},
  {8.9, 11.4, 12.4},
  {9.7, 11.5, 13.2},
  {9.8, 11.6, 13.1},
  {8.5, 10.3, 11.6},
  {7.6, 9, 11},
  {7.4, 8.8, 10.1},
  {7.1, 8.4, 9.5},
  {6.9, 8, 9},
  {6.4, 7.7, 8.6},
  {6.5, 7.8, 8.5},
  {6.4, 8.1, 8.2},
  {6.3, 7.8, 7.9},
  {6, 7.7, 7.6},
  {5.7, 7.5, 7.5},
  {4.4, 7.4, 7.2},
  {4, 7.2, 7},
  {3.3, 7.2, 6.9},
  {4.8, 7.7, 7.2},
  {7.3, 8.2, 8.5},
  {9, 8.9, 10.4},
  {10.1, 10.2, 12.4},
  {10.8, 11.8, 14},
  {11.6, 13, 15},
  {11.5, 13.7, 15.3},
  {11.8, 14.2, 15.3},
  {9.9, 13.6, 14.4},
  {9, 11.8, 12.7},
  {8, 10, 11.3},
  {7.5, 9.3, 10.7},
  {6.9, 9, 10.1},
  {6.7, 9, 9.5},
  {6.6, 8.9, 8.7},
  {6.7, 8, 8.2},
  {6.7, 7.8, 8},
  {6.6, 7.6, 8},
  {6.7, 8.1, 8},
  {6.4, 8.2, 8},
  {6.3, 7.9, 8},
  {6.2, 7.7, 7.9},
  {6.2, 7.5, 7.7},
  {6.1, 7.4, 7.4},
  {6.1, 7.2, 7.5},
  {6.1, 7.6, 7.7},
  {6.4, 7.7, 7.9},
  {7.1, 8.2, 8.3},
  {7.3, 8.1, 9.2},
  {7.6, 9, 10.4},
  {7.6, 10.1, 11.7},
  {8.6, 10.5, 12.7},
  {9, 11.5, 13.5},
  {9.8, 12, 13.7},
  {9.3, 11, 13.3},
  {8.7, 9.8, 12.4},
  {7.8, 9.3, 11.1},
  {7.9, 9.2, 9.5},
  {7.4, 9.1, 8.8},
  {6.9, 9.2, 8.6},
  {7.5, 8.9, 8.2},
  {7.4, 8.7, 8.1},
  {7.3, 8.9, 8},
  {6.6, 8.9, 8},
  {6.1, 8.1, 7.7},
  {5.8, 8, 7.5},
  {5.2, 7.7, 7},
  {6.1, 8.1, 6.6},
  {6.8, 8.7, 7.1},
  {7.6, 9, 8},
  {8.4, 9.5, 9.3},
  {8.4, 9.6, 10.9},
  {8.8, 10.9, 12.3},
  {9, 11.3, 13.5},
  {9.3, 11.4, 13.1},
  {9.6, 11.8, 13.3},
  {9.3, 12, 12.2},
  {9.4, 11.1, 13.1},
  {8.9, 10.8, 12.5},
  {8.4, 10.2, 11.8},
  {7.8, 9.8, 11},
  {7.5, 9.6, 10.2},
  {7.3, 9.4, 9.3},
  {7.1, 9.3, 8.8},
  {6.7, 9.1, 8.5},
  {6.9, 8.3, 8.4},
  {6.9, 8.1, 8.2},
  {6.8, 7.9, 8.2},
  {6.6, 7.5, 8},
  {6.5, 7.3, 7.9},
  {6.5, 7.5, 7.7},
  {6.5, 7.7, 7.6},
  {7.1, 8, 7.8},
  {7.3, 8, 8.2},
  {7.7, 8.4, 8.8},
  {8.4, 9.7, 9.4},
  {9.8, 11.1, 11},
  {10.6, 12.6, 13.3},
  {10.4, 13.7, 14.1},
  {11, 14.2, 15.6},
  {11.1, 14.2, 15.8},
  {10.3, 14.3, 14.3},
  {9.4, 12.9, 13.5},
  {7.7, 11.3, 11.7},
  {7.9, 9.9, 9.6},
  {7.7, 9.4, 8.1},
  {7.6, 8.7, 7.3},
  {7.4, 7.6, 7.2},
  {7.2, 6.6, 6.9},
  {6, 6.2, 5.8},
  {5.3, 6.4, 5.1},
  {4.9, 7.1, 4},
  {5.6, 7.1, 3.7},
  {4.7, 6, 3.1},
  {4.4, 5.7, 2.5},
  {4.7, 5.6, 3.3},
  {5.8, 5.5, 4.6},
  {9.1, 6.6, 5.4},
  {10.5, 9.3, 7},
  {12.8, 13.4, 12.2},
  {14.2, 15.7, 17.1},
  {15, 17.6, 19.4},
  {14.4, 17.6, 18.9},
  {13.2, 16.3, 16.9},
  {12.2, 15.7, 16.7},
  {12.8, 15.3, 17.7},
  {12.8, 14.7, 16.9},
  {10.7, 13.3, 15.1},
  {9.9, 12.8, 13.3},
  {10.3, 12.1, 11.9},
  {10.6, 10.9, 10.3},
  {9.5, 9.9, 9},
  {8.8, 9.7, 8.3},
  {8.9, 8.9, 7.9},
  {8.2, 8.4, 7.8},
  {7.4, 8.2, 7.3},
  {6.9, 8, 6.9},
  {6.6, 8, 6.8},
  {7.5, 7.5, 6.9},
  {7.5, 7.6, 7.2},
  {8.8, 8.3, 7.9},
  {9.6, 9.1, 9.6},
  {10.2, 9.5, 11.8},
  {10.2, 11.4, 13.9},
  {10, 12.4, 12},
  {10.2, 9.9, 12.3},
  {8.8, 8.5, 13.1},
  {8.5, 8.6, 12.9},
  {8.9, 8.5, 11.6},
  {8.6, 8.8, 12.3},
  {8, 8.9, 12.2},
  {7.4, 7.7, 11.4},
  {6.9, 7.3, 10.8},
  {6.6, 7.2, 10.1},
  {6.4, 6.9, 9.3},
  {6.5, 6.2, 8.6},
  {6.7, 5.9, 7.7},
  {7.3, 6, 7.3},
  {7.1, 5.7, 7.2},
  {6.7, 5.4, 6.8},
  {5.3, 5.4, 6.7},
  {5.7, 5.6, 5.7},
  {5.7, 5.7, 4.8},
  {5, 5.7, 5},
  {6.4, 6, 5.3},
  {7.8, 7.2, 5.7},
  {8.2, 8.8, 7.4},
  {9.6, 10.3, 9.7},
  {10.3, 12.3, 12.2},
  {11.8, 12.6, 15.6},
  {11.5, 13, 16.6},
  {12.1, 14.5, 15.8},
  {11.1, 14, 15.2},
  {10.5, 10, 15.1},
  {10.3, 8.4, 14.4},
  {9.8, 8, 13.1},
  {8.3, 7.5, 10.5},
  {7, 7.4, 9.8},
  {6.8, 7.4, 9.4},
  {7, 7.1, 9},
  {6.6, 6.8, 8.5},
  {6.6, 5.8, 8},
  {6.5, 5.4, 7.4},
  {6.2, 5.6, 7.3},
  {6.3, 6, 7.3},
  {5.6, 6.1, 7.4},
  {5.3, 5.9, 7.4},
  {6.4, 5.9, 7.5},
  {7.5, 6.9, 7.7},
  {7.7, 7, 8.1},
  {8.1, 8.3, 9.3},
  {8.9, 11, 10.9},
  {9.2, 11.6, 12.7},
  {9.2, 13.3, 13.2},
  {9.4, 11.2, 14.8},
  {9.1, 10.7, 12.7},
  {6, 9.8, 12.2},
  {6.1, 9.6, 11.2},
  {6.4, 8.9, 10.7},
  {6, 7.2, 10.6},
  {5.6, 6.6, 9.8},
  {5.4, 6.4, 9.1},
  {5.5, 5.9, 8.8},
  {5.6, 5.9, 8.4},
  {5.7, 5.8, 8},
  {5.5, 5.6, 7.7},
  {5.3, 5.6, 7.5},
  {5, 5.5, 7.1},
  {5.1, 5.6, 6.6},
  {4.9, 5.5, 6.5},
  {4.8, 4.6, 6.6},
  {4.6, 5.1, 6.6},
  {4, 6.2, 6.9},
  {4.9, 7.3, 7.8},
  {5.3, 8.3, 8.5},
  {6.5, 9.2, 10.9},
  {8.1, 10.5, 12.1},
  {8.6, 11.5, 12.2},
  {8.5, 12.1, 12.5},
  {8.4, 12.3, 12.5},
  {8.4, 11.8, 12.3},
  {8.2, 10.9, 11.9},
  {7.4, 9.6, 11.3},
  {6.7, 8, 10.5},
  {6.5, 7.1, 10.1},
  {6.1, 7.4, 9.9},
  {5.6, 7.5, 9.5},
  {5.3, 7.2, 9.5},
  {4.6, 6.7, 9.4},
  {4.1, 6.3, 9.3},
  {3.4, 5.7, 8.6},
  {2, 4.6, 7.5},
  {0.9, 2.9, 6.1},
  {0.7, 2.1, 4.7},
  {0, 2, 3.2},
  {1.3, 2.1, 3.3},
  {2.6, 3, 4.5},
  {5.1, 4.5, 6.7},
  {6.3, 7, 8.7},
  {7.2, 8.1, 10.8},
  {8.1, 10, 12.7},
  {9, 11.8, 12.7},
  {9.9, 12.6, 13.3},
  {10.5, 12.6, 13.4},
  {10.3, 12.2, 12.3},
  {10.1, 11.6, 12.2},
  {8, 10.3, 11.6},
  {5.1, 8.2, 10.4},
  {3.9, 7.3, 7.7},
  {3.3, 6.9, 5.9},
  {1.8, 5.5, 4.2},
  {1, 4.3, 3.1},
  {1, 4.6, 2},
  {0.9, 3.6, 1.2},
  {1.5, 3.1, 0.6},
  {1.5, 2.2, 0},
  {1.2, 1.6, -0.4},
  {0.6, 1.3, -0.9},
  {0.2, 0.8, -1.3},
  {0.3, 0.9, -1.6},
  {2.1, 1.6, -1.2},
  {5.8, 3.3, 1.4},
  {7, 6.4, 5.8},
  {7.9, 8.3, 9.5},
  {8.9, 10.3, 12.5},
  {10.1, 12, 14.9},
  {10.8, 13.4, 15.3},
  {11.4, 14, 15.3},
  {11.3, 13.9, 14.3},
  {10.1, 13, 12.9},
  {8.7, 10.8, 12.5},
  {7.2, 9.2, 11.4},
  {5.7, 8, 9.1},
  {4.7, 7, 6.6},
  {4.6, 6.1, 4.7},
  {3.5, 5.3, 3.4},
  {2.1, 4.5, 2.2},
  {1.7, 4.3, 1.4},
  {0.6, 3.5, 0.7},
  {0.7, 2.7, 0.1},
  {0.6, 2.1, -0.3},
  {0.3, 2.1, -0.7},
  {0.7, 2.2, -1},
  {0.8, 2.4, -1.4},
  {2.8, 2.6, -0.9},
  {6.6, 4.3, 3.2},
  {7.8, 6.9, 6.9},
  {9.1, 8.7, 10.3},
  {10.1, 11, 13.2},
  {11.3, 12.8, 14.7},
  {11.7, 14, 14.6},
  {11.6, 14.1, 14},
  {11, 13.6, 13.7},
  {10.3, 12.6, 13.6},
  {8.6, 11.6, 13},
  {6.8, 9.8, 11.5},
  {5, 8.7, 8.9},
  {5.9, 7.9, 6.5},
  {5.3, 7.6, 4.9},
  {2.8, 6.8, 3.3},
  {2.3, 5.1, 2.3},
  {1.8, 4.5, 1.3},
  {0.9, 3.8, 0.6},
  {0.8, 3.3, 0},
  {0.6, 2.3, -0.4},
  {0.8, 1.9, -0.9},
  {0.6, 2, -1.3},
  {0.9, 2.3, -1.4},
  {3.4, 3.2, -0.6},
  {6.9, 4.2, 3},
  {7.8, 6.8, 6.9},
  {8.9, 8.3, 11},
  {9.9, 10.6, 13.6},
  {10.7, 12.8, 14.6},
  {11.4, 13.5, 14.2},
  {11.7, 13.7, 14.4},
  {10.8, 12.9, 13.8},
  {10.4, 11.9, 13.7},
  {9.6, 11.4, 13.5},
  {8, 9.9, 11.8},
  {7.3, 8.9, 9.8},
  {6.6, 8.5, 7.5},
  {6.8, 7.7, 6},
  {6.4, 7.2, 5.2},
  {4.2, 6, 3.9},
  {3, 5.6, 3.1},
  {2.3, 5.1, 2.6},
  {2.2, 4.3, 1.6},
  {1.8, 3.8, 1.2},
  {2.2, 3.4, 0.7},
  {2, 3.7, 0.3},
  {2.5, 3.8, 0.2},
  {5, 4.6, 1.1},
  {7.5, 6.3, 4.4},
  {8.5, 7.3, 8.2},
  {9.4, 9.8, 11.6},
  {10.7, 11.7, 14.2},
  {12.3, 13.9, 15.8},
  {13.4, 14.7, 15.5},
  {13.2, 14.5, 15.4},
  {13.2, 14.4, 15.7},
  {13.3, 14, 15.4},
  {11.4, 12.9, 14.4},
  {8.9, 11.3, 12.8},
  {8.4, 10.1, 10.5},
  {8, 9.1, 8.7},
  {7.7, 8.5, 6.9},
  {7.4, 7.5, 5.7},
  {7.2, 7.8, 4.7},
  {6.9, 7.2, 4},
  {6.1, 7.3, 3.5},
  {5, 6.3, 3.3},
  {4.4, 5.8, 2.7},
  {4.2, 5.3, 2.6},
  {4.3, 5, 2.4},
  {5.3, 5.6, 2.8},
  {6.1, 6.7, 3.8},
  {7.1, 7.3, 5.8},
  {7.5, 8.2, 7.9},
  {8.3, 8.9, 10.3},
  {9.7, 10.7, 12.6},
  {10.4, 11.5, 14},
  {10.1, 11.6, 13.4},
  {8.5, 11, 13},
  {8.9, 10.5, 13},
  {9.1, 10.2, 12.8},
  {8.7, 10.1, 12.6},
  {8.2, 9.7, 11},
  {7.9, 9.7, 10.9},
  {7.2, 9.3, 9.7},
  {6.5, 9, 8.8},
  {6.1, 8.8, 8.3},
  {6.4, 8.4, 8.1},
  {6.6, 8.2, 8},
  {6.1, 8.3, 8},
  {5.7, 8.1, 7.6},
  {5.5, 7.9, 7.4},
  {5.7, 7.4, 7.1},
  {5.8, 7.7, 7},
  {5.6, 7.1, 6.9},
  {5.9, 7.1, 7.2},
  {6.1, 7.7, 7.6},
  {6, 7.9, 8.2},
  {6.3, 7.6, 9.5},
  {6.7, 7.5, 10.5},
  {6.8, 7.2, 10},
  {6.7, 7.1, 9.8},
  {6.7, 7.3, 9.4},
  {6.4, 7.4, 9.2},
  {5.5, 7.5, 8.5},
  {4.8, 6.7, 8},
  {4.2, 6.1, 7.1},
  {3.6, 5.5, 6.3},
  {3.4, 4.9, 5.9},
  {2.9, 4.6, 5.2},
  {2.3, 4.1, 4.7},
  {2.1, 2.8, 3.8},
  {2.1, 2.3, 2.9},
  {1.9, 2.3, 2.7},
  {2, 1.9, 2.6},
  {2, 2.1, 2.7},
  {2, 2.2, 2.8},
  {2, 2.2, 2.9},
  {2.2, 2.3, 3},
  {3, 3, 3.3},
  {3.5, 3.4, 3.9},
  {3.8, 4.1, 4.9},
  {3.9, 4.5, 5.7},
  {4.2, 5, 6},
  {4.8, 5.3, 6.8},
  {5, 6.4, 8.3},
  {5.6, 6.8, 9.4},
  {5.2, 6.9, 9.9},
  {5.7, 7, 10.3},
  {5.3, 6.7, 10.1},
  {4.6, 6.4, 9.4},
  {3.9, 5.5, 8.8},
  {3.9, 5, 7.8},
  {3.8, 5.3, 7.4},
  {4.3, 5.5, 6.4},
  {5.2, 6.2, 6.2},
  {5.5, 6.2, 5.9},
  {4.3, 6, 6},
  {4.2, 5.9, 4.9},
  {4.3, 5.8, 4.7},
  {4.5, 5.7, 5.1},
  {4, 5.3, 6.1},
  {4.3, 5.4, 6.7},
  {4.8, 5.8, 8.4},
  {4.7, 6.1, 9.1},
  {5.4, 6.7, 10},
  {5.8, 7.3, 10.3},
  {6.5, 7.9, 10.8},
  {6.7, 8.8, 11.3},
  {7.2, 9.3, 11.8},
  {7.5, 9.4, 12.2},
  {7.5, 9.4, 12.3},
  {7.6, 9, 12.3},
  {7.1, 8.3, 12.1},
  {6.6, 7.8, 11.8},
  {6.1, 7.6, 11.7},
  {5.8, 7.2, 11.2},
  {5.4, 6.9, 11.3},
  {5.2, 6.8, 11},
  {4.9, 6.7, 10.5},
  {3.5, 6.8, 9.8},
  {2, 6.6, 8.6},
  {1.6, 6.4, 8.2},
  {2, 6.2, 7.6},
  {1.8, 6, 6.9},
  {1.9, 5.9, 6.6},
  {2.4, 6, 6.3},
  {2.8, 5.9, 6.1},
  {3.5, 5.8, 6.3},
  {4.3, 5.9, 6.7},
  {5.3, 6.1, 6.9},
  {5.9, 6.7, 7.3},
  {6.7, 7.8, 7.7},
  {7.4, 8.8, 8.3},
  {7.8, 9.5, 9.1},
  {7.6, 9.8, 9},
  {7.8, 9.6, 9.3},
  {7.7, 9.5, 9.5},
  {7.3, 8.9, 9.4},
  {6.1, 8.5, 8.7},
  {6.2, 8, 8.2},
  {6.2, 7.9, 7.8},
  {5.9, 7.8, 7.5},
  {5.4, 7.4, 7.2},
  {5.4, 7.1, 7},
  {5.1, 7, 6.7},
  {4.9, 6.7, 6.6},
  {4.6, 6.8, 6.4},
  {4.6, 6.5, 6.4},
  {4.5, 6.5, 6.3},
  {4.8, 6.6, 6.1},
  {5, 6.8, 6.9},
  {5.2, 8.1, 8.2},
  {5, 8.4, 8.6},
  {5.1, 8.6, 10.2},
  {4.6, 8.7, 10.1},
  {4.5, 7.3, 8.5},
  {4.6, 6.6, 7.7},
  {4.7, 6.3, 7.6},
  {5.4, 8.2, 7.8},
  {5.2, 7.7, 7.9},
  {4.9, 6.7, 8.2},
  {4.1, 6.1, 8.2},
  {3.4, 5.3, 7.7},
  {2.7, 4.9, 7.2},
  {2.8, 4.6, 7},
  {3, 4.3, 6.8},
  {2.8, 4, 6.7},
  {3, 5, 6.5},
  {2, 5, 6.5},
  {2.2, 4.9, 6.5},
  {2.5, 4.9, 6.4},
  {3.3, 4.8, 6.5},
  {4, 4.7, 6.3},
  {4.6, 4.7, 6.2},
  {5.1, 4.9, 6.5},
  {5.9, 6.4, 7.3},
  {7.1, 8, 9.5},
  {9, 9.8, 11.8},
  {10.7, 11.7, 14},
  {11.6, 14.1, 16.2},
  {12.7, 15.8, 17.9},
  {13.1, 15.9, 16.7},
  {13, 16.2, 15.6},
  {12, 14.4, 15.7},
  {10.7, 13.3, 15.1},
  {9.4, 11.9, 13.5},
  {7.7, 10.8, 11.8},
  {6.8, 9.9, 9.9},
  {6.2, 9.3, 8.2},
  {6.4, 8.7, 7.6},
  {5.5, 8.1, 7},
  {5.8, 7.9, 6.1},
  {5.6, 8.1, 5.2},
  {5.2, 8.1, 4.8},
  {4.5, 7.2, 4.2},
  {4.9, 6.9, 3.9},
  {4.7, 6.1, 3.8},
  {6.2, 6.4, 4.3},
  {8.5, 7.5, 5.8},
  {10.4, 8.9, 7.4},
  {11.2, 10.6, 10.5},
  {12.1, 12.8, 14.4},
  {13, 14.7, 16.7},
  {13.6, 16, 16.6},
  {13.5, 16.6, 16.8},
  {12.1, 15.6, 15.8},
  {11.8, 14, 16.1},
  {11.6, 14.1, 16.9},
  {11.2, 13.9, 16.3},
  {10.7, 13.1, 15.5},
  {9.9, 11.9, 13.6},
  {8.9, 10.8, 10.3},
  {7, 10.3, 8.8},
  {6.5, 9.9, 7.8},
  {5.8, 9.7, 6.4},
  {5.5, 9.1, 5.5},
  {5.3, 7.8, 5.1},
  {5.3, 7.1, 4.2},
  {5.4, 6.7, 4.1},
  {4.8, 6.5, 3.7},
  {4.5, 7, 3.4},
  {5.3, 7.5, 3.2},
  {7, 8.1, 4.9},
  {9.2, 9.6, 6.8},
  {9.9, 11.4, 10.8},
  {11.2, 13.5, 13.9},
  {11.9, 14.4, 15.2},
  {12.7, 14.6, 15.5},
  {11.3, 14.1, 15.8},
  {9.7, 14.2, 14.7},
  {9.8, 13.8, 14.4},
  {9.6, 13.2, 13.7},
  {10, 12.7, 14},
  {9.7, 11.7, 13.4},
  {7.9, 10.5, 10.9},
  {6.4, 10.1, 9},
  {6.3, 10.1, 7.9},
  {7.1, 10, 7},
  {6.4, 9.7, 6.8},
  {5.7, 9.1, 6.3},
  {6.3, 8, 5.4},
  {7.5, 8.1, 5.3},
  {7.4, 7.7, 5.2},
  {7.6, 6.7, 5.3},
  {7.8, 7.2, 5.8},
  {7.9, 7.3, 6.1},
  {8.1, 8.2, 6.6},
  {8.8, 8.8, 7.1},
  {8.5, 8.9, 7.7},
  {7, 8.3, 7.8},
  {6, 7.5, 7.8},
  {5.7, 7.3, 8.1},
  {5.3, 6.8, 8.2},
  {4.7, 6.1, 8.2},
  {1.7, 5.6, 7},
  {1.6, 3.8, 5.4},
  {2.6, 3.7, 6},
  {2.5, 3.1, 5.8},
  {2.6, 3.2, 5.5},
  {2.6, 3.1, 5.2},
  {2.3, 3, 5},
  {1.9, 2.7, 4.5},
  {2.3, 1.7, 3.6},
  {1.7, 1.5, 3.4},
  {1.4, 1.3, 3.6},
  {0.4, 0.9, 3.6},
  {0, 0.5, 3.4},
  {0.2, 0.4, 3.2},
  {0.5, 0.3, 3},
  {1.5, 1, 3.4},
  {3.1, 2.1, 4},
  {3.5, 3.1, 5},
  {4.7, 4.1, 6.6},
  {6.1, 6.6, 7.8},
  {6.4, 8.2, 9.5},
  {7.1, 8.8, 11},
  {7.9, 10.4, 11.9},
  {8, 10.4, 12.7},
  {5.7, 9.2, 12.3},
  {6.5, 9.7, 8.9},
  {5.9, 9.2, 9},
  {4.5, 7.5, 8.3},
  {2.4, 5.7, 6.8},
  {2.4, 5.4, 5.4},
  {3.2, 5.1, 4.7},
  {2.9, 4.8, 3.9},
  {2.1, 4.1, 3.3},
  {2.7, 4.2, 3},
  {3.1, 4.2, 3.2},
  {3.3, 3.9, 2.9},
  {2.8, 3.5, 2.3},
  {2, 3, 1.7},
  {2.3, 2.7, 1.2},
  {2.3, 3.4, 1.1},
  {5.8, 4.2, 1.9},
  {7.5, 6.6, 5.4},
  {8.4, 9.1, 9.3},
  {10.2, 10, 12.4},
  {11.7, 12.1, 14.9},
  {12.5, 14.2, 17.3},
  {13.3, 14.8, 17.8},
  {12.9, 14.8, 16.6},
  {12.9, 14.8, 15.6},
  {11.8, 13.8, 15.4},
  {10.4, 12.4, 14.8},
  {9.7, 12.1, 14.4},
  {9.7, 11.5, 13.2},
  {9.5, 11.3, 11.7},
  {8.5, 10.7, 10.6},
  {7.8, 10.3, 9.3},
  {8.2, 9.8, 8.8},
  {7.8, 9.2, 8.7},
  {7.5, 8.9, 8.6},
  {8.2, 8.6, 8.5},
  {7.5, 8.3, 8.3},
  {6.6, 7.4, 8.1},
  {6.7, 7.1, 8.1},
  {7, 7, 8.1},
  {7.9, 7.2, 8.7},
  {8.9, 8.2, 10.2},
  {9.7, 8.9, 12.1},
  {10, 9.9, 13.4},
  {10.4, 11.1, 14.5},
  {10.4, 12, 13.7},
  {7.7, 12.4, 13.4},
  {5.8, 9.6, 10.1},
  {5.4, 8.2, 8.8},
  {5.4, 7.2, 8.8},
  {5.2, 6.8, 8.4},
  {5.2, 6.3, 8.2},
  {5.2, 5.9, 8.3},
  {5.2, 5.7, 8.1},
  {4.4, 5.6, 8},
  {4.4, 5.5, 7.8},
  {4.5, 5.3, 7.6},
  {4.5, 5.1, 7.6},
  {4.3, 4.8, 7.4},
  {4.3, 4.6, 7.3},
  {4, 3.9, 6.6},
  {3.7, 3.7, 6.5},
  {3.9, 3.8, 6.1},
  {4.1, 4.2, 6},
  {4.3, 5.3, 6.2},
  {5.1, 6.2, 6.9},
  {6, 6.7, 8},
  {6.7, 8.6, 9.7},
  {7.1, 9.3, 11.4},
  {7.8, 10.2, 13.1},
  {7.6, 11.1, 13.1},
  {7.2, 10.1, 11},
  {6.8, 9.8, 9.7},
  {6.4, 8.9, 10.3},
  {5.7, 8.4, 9.7},
  {5.3, 7.7, 9.3},
  {4.4, 6.8, 8.7},
  {4.1, 6.1, 8},
  {3.8, 5.6, 7.3},
  {3.3, 5.2, 7.1},
  {2.5, 4.4, 6.7},
  {2.2, 3.6, 6.5},
  {2.8, 3.5, 6.3},
  {2.7, 4, 6.5},
  {2.6, 4.4, 6.5},
  {2.6, 4.1, 6.2},
  {3, 4, 5.9},
  {3.4, 3.7, 5.8},
  {6.3, 4.8, 6},
  {7.8, 8.1, 8.7},
  {8.9, 10.2, 11.1},
  {10.1, 11.8, 13.7},
  {10.5, 13.2, 15.2},
  {11.1, 13.4, 16.2},
  {11.2, 13.7, 15},
  {10.6, 14, 14.7},
  {10.9, 13.9, 15.9},
  {9.7, 13.5, 15.7},
  {8.8, 12.2, 14.5},
  {7.2, 10, 12.9},
  {5.5, 8.1, 12.2},
  {4.6, 7, 12.3},
  {4.2, 6.3, 11.5},
  {3.8, 5.4, 10.7},
  {3.8, 4.8, 9.6},
  {3.8, 4.2, 7.4},
  {3.4, 3.4, 6.5},
  {2.8, 2.7, 5.8},
  {3.2, 2.1, 4.8},
  {3.1, 2, 3.9},
  {2.8, 1.7, 4.4},
  {2.6, 2.4, 4.6},
  {2.5, 3.3, 5.2},
  {2.8, 4.8, 6.6},
  {3.2, 6.4, 8},
  {4.1, 7.8, 8.9},
  {6, 9.1, 10.4},
  {6.6, 10.1, 11.7},
  {7.4, 11, 12.2},
  {8.3, 11.1, 12.1},
  {8.7, 11.1, 11.7},
  {8.2, 10.8, 11.8},
  {7.6, 10, 11.4},
  {5.9, 8.4, 10.3},
  {4.7, 6.8, 9},
  {3.7, 6.1, 7.3},
  {2.8, 5.1, 5.5},
  {3.2, 4.5, 4.4},
  {2.4, 4, 3.4},
  {2.5, 3.3, 2.7},
  {2.6, 3.3, 2.1},
  {3.5, 3.1, 1.8},
  {3.5, 3, 2.3},
  {3.7, 3.6, 3.2},
  {3.6, 3.7, 3.7},
  {3.7, 4.3, 4.2},
  {4.1, 4.7, 5},
  {4.7, 5.8, 6.3},
  {5.9, 6.8, 8.3},
  {6.1, 8.8, 9.7},
  {6.5, 9.6, 10.7},
  {7.7, 10.6, 11.2},
  {8, 11.3, 11.6},
  {8.4, 10.8, 12.2},
  {7.5, 11.1, 12.2},
  {7.3, 10.2, 11.9},
  {7.2, 9.4, 11.4},
  {6.9, 8.7, 10.8},
  {6.6, 8, 10.3},
  {6.3, 8, 10.2},
  {5.8, 7.9, 9.8},
  {5.5, 7.8, 9},
  {4.8, 7.6, 8.5},
  {3.9, 7.7, 7.9},
  {3.6, 7.6, 7.3},
  {4.9, 7.1, 7},
  {5.3, 7, 6.7},
  {5.4, 6.8, 6},
  {5.7, 6.3, 6},
  {6.1, 6.9, 6},
  {6.3, 7.8, 7.2},
  {6.6, 8.4, 9},
  {6.3, 8.7, 10.1},
  {6.5, 8.5, 10.6},
  {6.2, 8, 10},
  {5.7, 7.5, 9.3},
  {6, 7.7, 9.2},
  {6.3, 7.9, 9.7},
  {6.5, 7.9, 9.8},
  {6.4, 7.8, 9.8},
  {6.1, 7.4, 9.5},
  {6, 7.3, 9.2},
  {5.8, 7, 8.9},
  {5.5, 6.8, 8.5},
  {4.9, 6.3, 8.2},
  {4.2, 5.8, 8},
  {3.9, 5.2, 7.4},
  {3.8, 4.9, 6.9},
  {3.9, 4.9, 6.6},
  {3.9, 4.7, 6.5},
  {4.1, 4.7, 6.4},
  {3.9, 4.6, 6.2},
  {4, 4.6, 6.3},
  {4, 4.9, 6.4},
  {4.7, 5.3, 6.5},
  {5.1, 6.1, 6.9},
  {4.9, 5.8, 7.4},
  {5.5, 5.9, 8},
  {6.3, 6.6, 9.3},
  {7.4, 7.2, 11},
  {7.5, 7.7, 11.9},
  {8.9, 7.9, 11.8},
  {9.4, 8.9, 12.9},
  {8.1, 8.2, 12.5},
  {7.1, 7, 11.3},
  {6.5, 6.6, 10.3},
  {6.3, 6.6, 10},
  {6.3, 6, 9.7},
  {6.2, 5.4, 9.5},
  {5.7, 5.6, 9.3},
  {5.5, 5.6, 8.7},
  {5.3, 5.6, 8.4},
  {4.1, 5.5, 8},
  {3.7, 5.4, 7.8},
  {3.4, 4.7, 7.5},
  {3.2, 4.5, 7.3},
  {3.5, 4.2, 6.8},
  {5.4, 4.3, 6.5},
  {8.2, 5.4, 8.3},
  {8.9, 8.5, 10.1},
  {10.7, 12.2, 12.1},
  {12.4, 14.3, 15.2},
  {14.3, 15.8, 17.9},
  {15.6, 16.7, 19.3},
  {16.2, 18, 20.6},
  {16, 18.7, 20.5},
  {15.1, 19.1, 18.5},
  {14.9, 17.9, 18.5},
  {13.5, 16.5, 17.6},
  {12.4, 15.3, 17.1},
  {11.5, 13.6, 14.3},
  {10.9, 12.9, 11.8},
  {11.3, 12.3, 9.7},
  {10.9, 10.8, 8.3},
  {10.2, 10.1, 7.3},
  {8.9, 9.5, 6.6},
  {7.1, 8.4, 5.9},
  {6.7, 7.7, 5.4},
  {5.9, 7.5, 4.9},
  {6.1, 7.2, 4.3},
  {6.1, 7.2, 4},
  {8.5, 7.5, 4},
  {11.2, 8, 6.9},
  {12.5, 10.7, 10.8},
  {13.1, 13.1, 14},
  {14.2, 14.5, 17.1},
  {15.2, 16.7, 19.2},
  {16, 17.6, 19.5},
  {16.6, 18.1, 19.2},
  {16.1, 18, 19.5},
  {14.9, 17.9, 19.3},
  {14.9, 17.1, 19},
  {14, 16.7, 18.8},
  {13.1, 15.5, 17.6},
  {12.8, 14.1, 16.6},
  {12.5, 12.9, 14.1},
  {11.9, 12.3, 12.5},
  {11.8, 12.1, 10.9},
  {11.3, 10.9, 9.4},
  {9.8, 10.4, 8.6},
  {8.4, 9.9, 8},
  {7.5, 9.8, 7.3},
  {7.3, 9.6, 6.8},
  {7.1, 9.1, 6.2},
  {7.8, 8.8, 6},
  {9.8, 9.4, 6.2},
  {12, 10.7, 8.6},
  {12.3, 12.1, 11.5},
  {12.7, 13.2, 14.2},
  {13.4, 14.2, 17.1},
  {14.6, 14.5, 18.6},
  {14.6, 15.8, 18.4},
  {15.2, 16.9, 18.9},
  {15, 17.6, 19.2},
  {14.4, 17.2, 19.3},
  {15.1, 16.6, 18.8},
  {14.4, 16.2, 18.7},
  {13.4, 15.2, 17.5},
  {11.4, 13.9, 15.9},
  {10.3, 13.7, 14},
  {9.9, 13.3, 12.6},
  {9.6, 12.7, 11.5},
  {9.6, 12.6, 11.3},
  {9.5, 12.3, 11.2},
  {9.1, 12, 10.7},
  {9.3, 11.5, 9.8},
  {9.7, 11.2, 9.3},
  {9.1, 10.9, 8.6},
  {9.1, 11.1, 8.3},
  {10.6, 11.4, 8.9},
  {12.1, 12, 10.2},
  {12.9, 12.4, 11.9},
  {13, 13.1, 13.7},
  {13.2, 13.5, 15.2},
  {14.7, 14.5, 17.1},
  {15.6, 15.9, 19.8},
  {16.6, 17.4, 21.6},
  {17.1, 19.1, 22.2},
  {17.1, 20.4, 21.2},
  {15.3, 20.1, 20},
  {14.8, 18.5, 19.6},
  {13.6, 16.8, 18.4},
  {11.6, 14.8, 16.3},
  {10.5, 14.5, 14.3},
  {10.8, 13.4, 12.8},
  {10.1, 12.4, 11.7},
  {9.6, 11.9, 10.7},
  {9.4, 11.3, 9.9},
  {9.2, 10.9, 9.1},
  {8.9, 10.1, 8.4},
  {8.7, 9.7, 7.9},
  {8.6, 9.6, 7.5},
  {8.7, 9.4, 7.3},
  {11.7, 10.3, 8.2},
  {13.4, 10.8, 10.7},
  {14.1, 13.1, 14.7},
  {14.9, 15.3, 17.6},
  {15.8, 16.6, 19.8},
  {17.3, 18.3, 21.5},
  {18.3, 20.1, 22.1},
  {18.9, 21.9, 22.2},
  {19, 21.6, 22.9},
  {18.8, 21.3, 22.4},
  {17.7, 21, 22.2},
  {16.2, 19.9, 20.9},
  {15.1, 18.1, 19.3},
  {14.5, 16.5, 18},
  {13.5, 15.8, 15.7},
  {13.6, 15.1, 14},
  {13.4, 14, 12.8},
  {11.8, 13.7, 11.8},
  {10.1, 13.2, 10.8},
  {10, 12.5, 10.6},
  {9.8, 12.2, 11.1},
  {9.6, 11.4, 11.7},
  {10.6, 11, 11.9},
  {11.2, 11.4, 12.2},
  {12.4, 12.4, 12.6},
  {13.6, 13, 13.6},
  {14.6, 14.4, 14.9},
  {16.2, 16.2, 17.7},
  {17.5, 17.9, 20.4},
  {18.3, 19.3, 22.4},
  {19.5, 21.2, 23.9},
  {20.2, 22.6, 23.6},
  {20.7, 22.5, 23.6},
  {20.6, 21.9, 23.1},
  {19.9, 21.7, 22.7},
  {18.5, 20.6, 22.5},
  {16.7, 19.2, 21.3},
  {16.1, 17.7, 19.5},
  {15.7, 16.9, 17.3},
  {15.5, 15.9, 15.2},
  {14.9, 15.6, 14},
  {13.9, 15.1, 12.9},
  {12, 14.3, 11.9},
  {11.2, 13.5, 11.4},
  {11.5, 12.9, 10.8},
  {11, 12.3, 10.4},
  {10.6, 12.4, 9.7},
  {10.6, 12.5, 9.6},
  {12.7, 12.9, 9.8},
  {15.6, 13.8, 12.2},
  {16.4, 15.4, 15.4},
  {17.7, 17.2, 18.9},
  {18.7, 19.6, 21.8},
  {19.7, 21.1, 23.6},
  {19.8, 22.2, 23.6},
  {21.2, 22.1, 23.6},
  {_, 22, 23.7},
  {_, 22, 23.4},
  {_, 21.2, 22.9},
  {_, 20.9, 23.2},
  {_, 19.8, 21.9},
  {_, 18.4, 20.3},
  {_, 17.4, 17.8},
  {_, 17.5, 15.8},
  {_, 16.6, 14.5},
  {_, 15.6, 13.5},
  {_, 14.9, 12.8},
  {_, 14, 11.8},
  {_, 13.3, 11.4},
  {_, 13, 10.6},
  {_, 12.4, 10.3},
  {_, 12.6, 10.5},
  {_, 13.9, 11.1},
  {_, 15.1, 13.3},
  {_, 16, 15.7},
  {_, 17.9, 18.3},
  {_, 19.1, 21.1},
  {_, 19.7, 22.4},
  {19.3, 20.4, 22.9},
  {18.7, 20.8, 22.3},
  {18.6, 20, 22.8},
  {18, 20.8, 22.5},
  {17.4, 19.7, 21.5},
  {16.7, 18.7, 20.8},
  {16.2, 18.1, 20.5},
  {15.5, 16.8, 19.5},
  {14.6, 16, 17.5},
  {13.6, 15.5, 15.1},
  {14, 15.2, 14.4},
  {11.2, 12.1, 13.9},
  {10.2, 8.9, 13},
  {9.6, 9, 12.2},
  {7.6, 8.9, 11.1},
  {6.7, 8.5, 9.7},
  {6.4, 8.4, 8.5},
  {6.6, 9.1, 7.8},
  {8.9, 9.1, 8},
  {11.4, 9.6, 9.5},
  {12.2, 11.3, 12.3},
  {13.2, 13.7, 14.7},
  {14.7, 15.9, 17.8},
  {16.5, 18.2, 20.2},
  {17.9, 19.8, 21.9},
  {18.2, 20.6, 22.1},
  {17.3, 18.9, 19.7},
  {16.8, 17.2, 18.8},
  {15.8, 13.3, 16.2},
  {13.4, 12.1, 14.9},
  {12.7, 11.6, 13.2},
  {11.3, 10.8, 12.4},
  {9, 10.3, 11.9},
  {8.7, 9.8, 11},
  {8.7, 10, 9.9},
  {9.4, 9.7, 9.7},
  {9.3, 8.9, 9.7},
  {8.8, 8.5, 9.5},
  {8, 8.5, 9.3},
  {7.8, 8.3, 9},
  {7.6, 8.1, 8.8},
  {7.8, 8.2, 8.8},
  {8.7, 9.6, 9.3},
  {9.3, 10.3, 10.2},
  {9.7, 12.8, 11.1},
  {11.7, 14.1, 13.2},
  {12.7, 14.8, 15.8},
  {12.8, 16.5, 18},
  {12.5, 16.8, 17.4},
  {9.5, 17.6, 14},
  {9.9, 17, 13.7},
  {11.6, 17.4, 15.4},
  {11.2, 16, 15.2},
  {10.7, 13.6, 14.4},
  {9.1, 12.2, 13.5},
  {7.8, 10.8, 12.7},
  {6.9, 9.7, 10.6},
  {7.2, 9.2, 9.1},
  {7.6, 9.2, 8},
  {7.3, 9.1, 7.1},
  {6.6, 8.8, 6.3},
  {6.7, 8.6, 5.7},
  {6.2, 8.1, 5},
  {6, 8, 4.4},
  {6.5, 7.5, 3.8},
  {6.3, 7.7, 3.4},
  {9.4, 8.8, 4.2},
  {11.3, 10.8, 6.5},
  {11.8, 12.5, 10},
  {13, 12.9, 13.4},
  {13.9, 13.9, 15.2},
  {15.5, 16.1, 18.3},
  {15.9, 17.3, 20.1},
  {15.4, 17.6, 21},
  {14.3, 17.6, 19.8},
  {13.5, 17.4, 18.7},
  {14.4, 17.5, 18},
  {14, 16.3, 18.9},
  {12.3, 16.2, 18.4},
  {10.6, 14.6, 15},
  {10, 12.7, 11.9},
  {9.7, 11.8, 9.9},
  {8.7, 10.8, 8.4},
  {7.4, 9.9, 7},
  {7.2, 9.1, 5.7},
  {6.1, 9, 4.9},
  {5.2, 8.5, 4.3},
  {4.9, 8.1, 3.7},
  {4.8, 7.9, 3.1},
  {4.9, 7.3, 2.6},
  {8.9, 7.6, 3.4},
  {11.1, 9, 6.6},
  {11.8, 12, 10.9},
  {13.5, 14, 14.9},
  {14.3, 15, 17.8},
  {15.2, 16.4, 19.5},
  {15.4, 17.7, 19.8},
  {15.9, 18, 19.2},
  {15.5, 17.9, 19},
  {15.9, 18.1, 19.5},
  {15.4, 17.8, 19.5},
  {15.1, 16.9, 19},
  {14.7, 16, 18.6},
  {14.2, 14.3, 16.7},
  {13.7, 13.4, 14.1},
  {12.4, 12.9, 12},
  {11.8, 12.1, 10.3},
  {11.5, 11.4, 8.8},
  {11.2, 10.6, 7.4},
  {10.3, 10.4, 6.8},
  {8, 9.8, 6.1},
  {6.5, 9.6, 5.2},
  {5.2, 8.9, 4.8},
  {5.8, 8.5, 4.3},
  {9.3, 8.6, 5.6},
  {10.9, 9.2, 9.5},
  {11.4, 11.5, 12.9},
  {13.2, 13.1, 16.6},
  {13.8, 13.8, 16.9},
  {14.2, 14.6, 17.8},
  {14.7, 15.2, 18.4},
  {15.1, 15.7, 19.1},
  {15.5, 15.9, 19.7},
  {14.5, 16, 19.8},
  {13.8, 15.6, 19.2},
  {13.6, 15, 18.3},
  {12.6, 13.8, 16.9},
  {11.7, 12.5, 16.5},
  {10.6, 12.1, 15.2},
  {9, 11.2, 14.9},
  {9.5, 10.9, 14.1},
  {8.9, 10.6, 13.2},
  {8.4, 9.7, 12.7},
  {7.7, 8.4, 11.8},
  {7.4, 6, 11.5},
  {7.2, 4.9, 11.1},
  {6.8, 5, 10.4},
  {6.3, 5.2, 9.6},
  {7.2, 5.8, 10.1},
  {7.5, 6.2, 11.4},
  {8.2, 7.1, 12.2},
  {8.3, 7.8, 12},
  {8.4, 8.4, 11.9},
  {8.8, 9.5, 11.7},
  {8.1, 11.8, 13.2},
  {7.1, 11.5, 13},
  {6.5, 12.6, 12.6},
  {7.3, 13, 12.9},
  {8.2, 12.6, 14.2},
  {7.8, 12.1, 13.3},
  {7.4, 10.5, 11.9},
  {7.3, 9.3, 11.4},
  {7, 8.8, 11},
  {6.8, 8.1, 11},
  {6.8, 8.4, 11.1},
  {6.7, 8.1, 10.9},
  {6.6, 8.2, 10.5},
  {6.4, 8.2, 9.2},
  {6.3, 7.8, 8.3},
  {6.6, 7.3, 8.3},
  {6.6, 7.1, 8.3},
  {6.4, 6.9, 7.8},
  {6.4, 7, 8.2},
  {6.6, 8, 8.6},
  {6.4, 8.4, 8.9},
  {5.8, 8.4, 9.4},
  {6.1, 9.1, 10.4},
  {6.6, 9.7, 11.3},
  {8.1, 10, 11.6},
  {8.5, 10.9, 12},
  {9.4, 11.2, 12.8},
  {9.6, 11.1, 13.2},
  {9.3, 10.9, 13.2},
  {8, 10.6, 12.9},
  {7.9, 10, 12.4},
  {7.1, 9.2, 11.7},
  {7, 8.4, 11.1},
  {7.1, 7.9, 10.5},
  {6.8, 7.7, 9.7},
  {6.9, 7.5, 9.6},
  {6.9, 7.1, 9.2},
  {6.6, 7.3, 9},
  {5.8, 7.3, 8.6},
  {5.3, 7.1, 7.8},
  {4.8, 6.8, 7},
  {4.4, 6.2, 6.3},
  {7.4, 6.1, 6.6},
  {8.5, 7.1, 9.6},
  {9, 9.7, 12.5},
  {10.6, 11.8, 15.1},
  {12.1, 13.2, 16.6},
  {11.8, 14.6, 17.8},
  {11.8, 14.8, 15.5},
  {12.2, 15, 16.7},
  {11.3, 15.3, 16.5},
  {12, 14.6, 15.8},
  {11.7, 14.4, 15.7},
  {11.2, 13.7, 14.8},
  {10.4, 12.5, 14.5},
  {10, 10.7, 13.6},
  {9.6, 10.4, 12.8},
  {8.3, 10.2, 12.4},
  {8.5, 9.9, 11.6},
  {7.3, 10.1, 10.9},
  {7.1, 9.3, 10.5},
  {6.9, 9.2, 10},
  {7.1, 8.5, 9.6},
  {7.3, 8.4, 9.4},
  {7.2, 8.5, 9.2},
  {7, 7.9, 9.1},
  {8.5, 8.4, 9.1},
  {10.2, 9.7, 9.9},
  {10.9, 10.9, 12.5},
  {11.6, 11.7, 14.7},
  {12.2, 12.9, 16.3},
  {12.8, 15, 17.7},
  {13.4, 16.4, 17.6},
  {14.1, 16.6, 18},
  {14.2, 17.4, 18.2},
  {13.8, 17.4, 17.7},
  {13.3, 16.9, 17.1},
  {12.4, 15.2, 16.4},
  {11.2, 13.6, 15.9},
  {9.9, 12.3, 14.7},
  {8, 11.2, 13.5},
  {7.3, 10.7, 11.4},
  {6.6, 9.9, 9.8},
  {6.5, 9.1, 8.4},
  {6.1, 8.9, 7.3},
  {6.8, 8.1, 6.4},
  {7.8, 8.2, 6.6},
  {7.2, 8.4, 6.9},
  {7.3, 7.8, 7.1},
  {8, 8, 7.2},
  {8.9, 9.1, 7.6},
  {9.8, 9.8, 9.2},
  {11.1, 10.9, 11.7},
  {12.5, 13.2, 14.5},
  {13.4, 14.1, 17.6},
  {14.4, 16.2, 18.5},
  {15.3, 17.2, 18.8},
  {15.5, 18, 19.2},
  {16.1, 18.2, 19.9},
  {16.1, 18.4, 19.6},
  {15.2, 18, 19.4},
  {13.4, 16.6, 18.6},
  {12.9, 15, 17.4},
  {11.6, 14.2, 16.7},
  {9.3, 13.3, 14.5},
  {9.8, 12.7, 12.1},
  {9.4, 12, 10.3},
  {8.9, 11.6, 9.3},
  {9.9, 11.4, 9},
  {9.3, 10.9, 8.6},
  {9.3, 10.8, 8.9},
  {9.4, 11, 9.3},
  {9.6, 10.5, 9.3},
  {9.9, 10.2, 9.3},
  {10.6, 11, 9.8},
  {11.6, 11.9, 10.6},
  {12.1, 13, 12.2},
  {12.7, 13.3, 13.4},
  {13, 14, 14.1},
  {10.3, 14, 15},
  {9.3, 11.8, 12.6},
  {9.4, 11.3, 12.5},
  {9, 10.7, 12.5},
  {8.8, 10.2, 12.1},
  {9.3, 10.4, 12.1},
  {10, 11.1, 12.8},
  {10, 11.3, 12.6},
  {9.1, 9.8, 12.3},
  {8.8, 9.6, 11.5},
  {8.9, 9.5, 11.5},
  {8.9, 9.3, 11.5},
  {9, 9.4, 11.5},
  {9.1, 9.3, 11.4},
  {9, 8.7, 11.3},
  {8.7, 8.4, 11.1},
  {7.1, 8.2, 10.8},
  {6.3, 8.9, 10.5},
  {7.3, 9.4, 10.5},
  {9, 9.4, 10.9},
  {9.5, 10.1, 12},
  {11.4, 12, 14.2},
  {12.4, 13.3, 15.8},
  {13.4, 14.7, 17.8},
  {14.6, 17, 19.1},
  {15.1, 17.5, 17.4},
  {15.1, 17.1, 16.8},
  {13.9, 16.7, 16.8},
  {14.5, 15.9, 17.1},
  {13.6, 16, 17},
  {12.8, 15, 16.9},
  {12.4, 14.2, 16.4},
  {11.7, 13, 15.8},
  {11.2, 12.5, 14.6},
  {11.3, 12.8, 13.1},
  {11.2, 12.6, 12.1},
  {11.1, 12.5, 12.2},
  {10.6, 12.2, 12.3},
  {9.9, 12.3, 12.3},
  {8.8, 12, 12.1},
  {9.4, 11.3, 11.8},
  {10.1, 11.4, 11.5},
  {10.1, 11.6, 11.1},
  {10.5, 12.3, 11.6},
  {11.1, 12.8, 12.5},
  {12, 13.6, 14.2},
  {12.4, 14.2, 15.5},
  {13, 15.2, 16.1},
  {12.8, 15.4, 16.6},
  {13.6, 15.7, 17.8},
  {13.1, 15.7, 18.2},
  {13.5, 14.6, 18.1},
  {13.5, 15.6, 18.5},
  {13.6, 15.4, 18.2},
  {12, 15.2, 16.9},
  {11.3, 13.3, 13.2},
  {10.9, 11.9, 11.8},
  {9.1, 10, 11.1},
  {8.8, 9.5, 10.9},
  {8.4, 9.5, 10.8},
  {8.5, 9.1, 10.6},
  {8.7, 8.9, 10.1},
  {8, 8.4, 9.9},
  {7.7, 7.5, 9.7},
  {7.3, 7.1, 9.4},
  {7.1, 7.4, 9.3},
  {7.3, 8.1, 9.3},
  {9.4, 9, 10.1},
  {10.7, 9.5, 11.2},
  {11.2, 10.4, 12.5},
  {12.9, 12.1, 15.1},
  {14.3, 13.8, 16.4},
  {14.6, 15.9, 17.9},
  {14.3, 16.9, 17.5},
  {15.7, 17.1, 17.1},
  {13.4, 15.8, 16.3},
  {13.4, 13.6, 15.5},
  {13.3, 12.3, 14.4},
  {12.7, 11.6, 14.5},
  {11.9, 11.1, 13.9},
  {10.1, 10.9, 13.2},
  {9.5, 10.9, 11.8},
  {9.1, 10.3, 11.4},
  {8.9, 9.8, 11.3},
  {8.7, 9.7, 10.5},
  {8.6, 9.6, 10.1},
  {8.1, 9.4, 10},
  {7.7, 8.9, 9.8},
  {7.5, 8.5, 9.6},
  {7.6, 8.2, 9.5},
  {7.2, 8.3, 9.4},
  {6.8, 8.5, 9.4},
  {7, 8.4, 9.4},
  {7.4, 8.3, 9.4},
  {7.3, 8.4, 9.4},
  {7.1, 8.6, 9.5},
  {8.3, 9.8, 9.7},
  {10.5, 10.1, 10.6},
  {11.5, 10.3, 12.1},
  {10.7, 10, 13.4},
  {11.3, 10.2, 13.2},
  {10.8, 10.8, 13.4},
  {11, 10.6, 13.8},
  {10.5, 10.3, 13.7},
  {11.1, 10.4, 12.5},
  {11.2, 10.3, 11.7},
  {9.8, 10.1, 10.9},
  {9.8, 10, 10.1},
  {8.7, 10, 9.4},
  {7.7, 9.9, 8.8},
  {7.2, 9.6, 8.6},
  {6.7, 8.8, 7.5},
  {6.4, 8, 6.4},
  {5.5, 7.2, 5.6},
  {6.9, 7, 4.9},
  {9.4, 8.2, 5.5},
  {10.6, 9.1, 8.2},
  {10.9, 11.5, 11},
  {12.7, 13.4, 14.6},
  {13.7, 14.9, 17},
  {15, 16.6, 18.5},
  {16.1, 18.3, 20.2},
  {16.6, 19.4, 20.3},
  {16.4, 19.9, 20.2},
  {16.1, 20, 20},
  {14.7, 19.5, 20},
  {13.9, 18.2, 19.4},
  {13.1, 16.9, 18.6},
  {12.7, 14.9, 16.6},
  {12.3, 13.3, 14.3},
  {11.9, 12.2, 12.3},
  {11.1, 11.4, 10.8},
  {9.4, 10.5, 9.7},
  {8.1, 9.9, 8.9},
  {7.4, 9.1, 8.2},
  {6.9, 8.7, 7.5},
  {6.7, 8, 7},
  {6.6, 7.7, 6.6},
  {7.6, 7.5, 6.2},
  {10.8, 7.9, 7.2},
  {11.8, 9.1, 9.7},
  {12.8, 11.9, 12.8},
  {13.7, 14.2, 15.8},
  {15, 16.1, 18.4},
  {16, 17.7, 20.2},
  {17, 19.4, 20.1},
  {16.9, 19.7, 20.4},
  {17.3, 19.9, 20.9},
  {16.9, 18.9, 20.2},
  {16.5, 18.7, 20},
  {15.7, 18.2, 19.5},
  {14, 17.2, 18.8},
  {12.9, 15.5, 17.1},
  {11.8, 14.3, 15},
  {11.2, 13.3, 13.4},
  {10.6, 12.6, 12.3},
  {9.8, 12.1, 11.4},
  {9.4, 11.4, 10.5},
  {9.1, 10.9, 9.8},
  {8.9, 10.4, 9.2},
  {8.7, 10.5, 8.7},
  {8.5, 10.1, 8.3},
  {9.6, 10.2, 8},
  {12.9, 10.7, 8.8},
  {14.2, 12, 11.7},
  {14.7, 14.3, 14.9},
  {16, 16.1, 17.9},
  {17.3, 17.9, 20.8},
  {18.4, 19.6, 22.8},
  {19.6, 21.3, 22.1},
  {19.7, 21.4, 22.9},
  {20, 21.4, 22.8},
  {19.3, 21.2, 22.6},
  {19.6, 19.9, 22},
  {18.6, 18.9, 21.4},
  {16.5, 18.4, 20.5},
  {15.5, 17.6, 19.9},
  {14.8, 16, 17.8},
  {14.6, 15.5, 15.9},
  {14, 15.1, 14.7},
  {13.2, 14.8, 14},
  {12.9, 14.4, 13.4},
  {12, 14.1, 13},
  {11.3, 13.4, 12.3},
  {11.9, 13.6, 12},
  {11.7, 13.7, 12},
  {12.1, 14, 12.1},
  {13.8, 14.3, 12.9},
  {15.3, 15.4, 14.4},
  {16.2, 16.9, 17.3},
  {17.3, 18.1, 20.1},
  {17.9, 18.8, 21.4},
  {18, 20.2, 21.9},
  {19.4, 20.7, 22.3},
  {20.2, 22, 23.6},
  {19.7, 22.2, 23.2},
  {18.9, 21.7, 23},
  {18.8, 21.3, 22.7},
  {17.9, 20.3, 22},
  {17.1, 19.2, 21},
  {15.8, 16.9, 20},
  {14.3, 16.3, 17.2},
  {15, 16.6, 15.7},
  {14, 16.2, 14.3},
  {12.7, 15.5, 12.6},
  {12.4, 14.6, 12.3},
  {11.6, 14.8, 11.6},
  {12.5, 14.2, 11.6},
  {12.3, 13.5, 11.2},
  {12.4, 13.3, 11.1},
  {13.1, 13.3, 11.6},
  {14, 13.7, 11.9},
  {15, 13.4, 12.2},
  {15.2, 14.5, 13.2},
  {15.6, 14.4, 14.6},
  {15.8, 14.9, 16.5},
  {15.7, 15.5, 17.8},
  {15.8, 14.8, 17.5},
  {15.4, 15.1, 17.4},
  {15, 14.7, 17.9},
  {14.4, 14.7, 17.8},
  {13.8, 15, 16.6},
  {12.5, 14, 15.4},
  {10.9, 12.1, 13.5},
  {10.2, 11.5, 12.6},
  {10.1, 10.6, 12.4},
  {10.3, 9.2, 12.1},
  {9.7, 9, 11.9},
  {8.8, 9, 11.6},
  {7.9, 8.8, 10.7},
  {6.8, 8.6, 9.5},
  {6.2, 8.5, 8.6},
  {6.7, 8.4, 7.9},
  {7.7, 8.4, 7.3},
  {8.4, 9, 7.1},
  {9.6, 9.5, 8.3},
  {11.6, 10.1, 9.2},
  {12.5, 11.3, 10.8},
  {13.3, 13.9, 13.8},
  {14.8, 16.4, 17.4},
  {16.7, 18.1, 19.8},
  {18, 19.9, 21.8},
  {18.6, 19.7, 23.3},
  {19, 21.6, 23.6},
  {19.3, 22.1, 22.6},
  {18.7, 21.5, 21.9},
  {16.7, 20.5, 21.8},
  {15.6, 19.6, 20.9},
  {14.9, 17.6, 18.9},
  {14.2, 15.6, 16.3},
  {11.6, 13.9, 14.3},
  {11.2, 13.3, 12.8},
  {11.2, 12.6, 11.9},
  {11.1, 12.5, 11.1},
  {11.1, 12.1, 10.4},
  {11, 11.5, 9.8},
  {10.3, 10.9, 9.3},
  {10.2, 10.5, 8.8},
  {11.2, 10.7, 8.5},
  {14.5, 11.2, 9.3},
  {15.5, 12.5, 12.6},
  {15.3, 15.3, 15.9},
  {17.1, 17.2, 19},
  {18.3, 18.7, 21.6},
  {19.4, 20.6, 23.8},
  {20, 22.4, 23.6},
  {20.2, 23.3, 23.4},
  {20.4, 23.2, 24},
  {20.3, 23.2, 24.1},
  {20.3, 22.6, 24.4},
  {18.9, 21.8, 23.6},
  {16.9, 20.3, 22.1},
  {15.1, 18.7, 20.5},
  {13.7, 17.5, 18.4},
  {13.1, 16.6, 16.5},
  {12.9, 15.7, 15.1},
  {12.6, 15.4, 14.2},
  {12.3, 14.6, 13.4},
  {12, 14, 12.7},
  {11.7, 13.2, 12.2},
  {11.5, 12.9, 11.6},
  {11.6, 12.4, 11.2},
  {12.4, 12.7, 11.2},
  {15.2, 13.9, 12.3},
  {16.8, 15, 13.3},
  {17.5, 16.8, 14.7},
  {18.1, 18.7, 16.9},
  {18.5, 20, 20.7},
  {19.7, 21.8, 23.6},
  {20.2, 22.9, 24.5},
  {21.1, 23.5, 24.5},
  {21.2, 23.7, 24.7},
  {21.3, 23.7, 24.4},
  {21.5, 22.9, 24.3},
  {19.7, 22.4, 24},
  {17.8, 21.1, 22.7},
  {17.3, 19.5, 21.2},
  {15.3, 18.4, 20},
  {14.5, 17.9, 19.3},
  {14.8, 16.8, 18.5},
  {14.7, 16.3, 17.7},
  {14.9, 16.2, 17.1},
  {15.5, 15.2, 16},
  {15.9, 14.4, 14.8},
  {14.3, 14.1, 14.6},
  {13.3, 13.7, 13.8},
  {14, 13.9, 13.2},
  {17.5, 14.4, 14.5},
  {19, 15.4, 16.9},
  {19, 18.2, 20.2},
  {20.1, 19.9, 22.6},
  {21.1, 21.9, 24.9},
  {22.2, 23.5, 27},
  {23.1, 25.1, 26.9},
  {23.3, 25.9, 27.1},
  {23.6, 26, 27.2},
  {23.3, 25.8, 26.8},
  {22.6, 25.1, 26.2},
  {21, 24.1, 26.1},
  {19.7, 23, 25.1},
  {17.8, 21.4, 23.5},
  {16.2, 20.2, 21.3},
  {15.6, 19, 19.1},
  {14.8, 17.8, 18},
  {15, 17.4, 17.3},
  {15.2, 16.3, 16.3},
  {14.7, 15.4, 15.5},
  {14, 15.6, 14.7},
  {14.9, 15.6, 14.2},
  {14.1, 15.4, 13.8},
  {14.9, 15.2, 13.5},
  {18.2, 15.5, 14.4},
  {20.1, 17, 17.6},
  {20.2, 19.5, 20.9},
  {21.3, 20.8, 23.4},
  {22.5, 22.8, 26},
  {23.4, 24.7, 27.9},
  {24.3, 26.5, 28.6},
  {24.6, 26.9, 28.4},
  {24, 26.5, 28.7},
  {23.8, 24.9, 28.5},
  {22.8, 24.9, 28.1},
  {21.5, 23.4, 26.8},
  {20.7, 23.1, 25.5},
  {20.1, 21.4, 24},
  {17.2, 20.7, 21},
  {16.6, 19.4, 19},
  {16.2, 18.1, 17.5},
  {15.6, 17.4, 16.6},
  {15.9, 16.9, 15.7},
  {15.3, 16.2, 15.1},
  {15.6, 16.5, 14.8},
  {15, 16.5, 14.4},
  {15.4, 16.2, 13.7},
  {16.4, 15.9, 13.3},
  {19.3, 16.2, 14.4},
  {20.2, 17.6, 17.4},
  {20.4, 19.9, 20.7},
  {22.1, 21.4, 23.3},
  {23.5, 23.2, 26.1},
  {24.1, 25, 28.2},
  {24.8, 26.8, 29.1},
  {24.7, 27.3, 29.2},
  {23.6, 27.6, 29.3},
  {23.8, 27, 29.1},
  {23.6, 26.6, 28.9},
  {22.4, 25.9, 27.8},
  {20.8, 24.9, 26.7},
  {19.9, 23, 24.8},
  {17.5, 21, 21.9},
  {16.9, 20.8, 19.2},
  {16.6, 20.4, 17.8},
  {16, 18.9, 16.6},
  {15.7, 17.7, 15.8},
  {15.5, 16.7, 15},
  {15.1, 16.1, 14.3},
  {14.3, 15.6, 13.7},
  {14.5, 15.6, 13.2},
  {15.4, 15.9, 13},
  {18.7, 16.1, 14},
  {20.4, 17, 17.8},
  {20.9, 19.8, 20.6},
  {22.5, 21.6, 23.5},
  {23.5, 23.7, 26},
  {23.9, 25.3, 28.1},
  {24.2, 26.2, 28.3},
  {24.4, 26.7, 28.3},
  {24.1, 26.9, 28.5},
  {23.9, 26.6, 28.4},
  {22.7, 25.4, 27.4},
  {22.4, 24.5, 26.8},
  {21, 23.5, 26},
  {19.9, 22.1, 25.1},
  {19, 20.7, 22.9},
  {18.6, 20.4, 21},
  {18.3, 20.6, 19.8},
  {18.5, 20.1, 19.4},
  {17.7, 17.2, 19.2},
  {17.5, 14.1, 18.6},
  {16.3, 13.9, 19.5},
  {15.8, 13.8, 19.3},
  {13.9, 13.7, 18},
  {14.3, 13.9, 16.7},
  {16.1, 14.1, 17.2},
  {17.3, 14.8, 18.4},
  {17.8, 17, 20.3},
  {19, 18.4, 21.9},
  {20.2, 20, 23.9},
  {21.9, 21.7, 25.7},
  {22.1, 23.6, 27.1},
  {20.4, 23.9, 27.2},
  {20.2, 21.7, 24.2},
  {18.5, 19.6, 17.8},
  {16.7, 19, 17.4},
  {17, 18.6, 17.1},
  {16.6, 16.9, 17.9},
  {16.3, 15.3, 17.7},
  {15.9, 14.3, 17.5},
  {15.5, 14.4, 17.2},
  {15, 14.2, 17.1},
  {14.5, 14.2, 17.1},
  {13.7, 13.7, 17},
  {13.1, 12.7, 16.3},
  {12.4, 11.5, 15.7},
  {11.9, 10.5, 15.1},
  {11.4, 9.7, 14.5},
  {12.5, 9.7, 13.9},
  {13.2, 10.5, 13.8},
  {13.7, 11.5, 15.6},
  {14.3, 14.5, 16.7},
  {15.6, 16.9, 18.4},
  {17.2, 18.1, 20.6},
  {17.4, 19.3, 21.2},
  {17, 19.8, 20.9},
  {16, 20.1, 20.4},
  {15.6, 19.8, 20.6},
  {15.9, 19.3, 19.9},
  {15.7, 18.4, 19.7},
  {15.7, 17.7, 19.8},
  {15.2, 17.4, 19.6},
  {15, 15.8, 18.9},
  {14.9, 15, 18.3},
  {14.5, 15.7, 17.5},
  {14.1, 15.3, 16.6},
  {13.7, 15.2, 16.3},
  {13.2, 15.3, 16.1},
  {13, 14.9, 15.8},
  {12.8, 14.5, 15.6},
  {12.2, 13.7, 15.4},
  {11.8, 13.4, 15},
  {12.3, 13.8, 15.1},
  {13.2, 14.5, 15.4},
  {14.9, 15.3, 16.8},
  {16.1, 16.2, 18.9},
  {16.8, 17.9, 20.5},
  {17.8, 19.2, 21.9},
  {18, 20.2, 21.7},
  {17.9, 20.7, 21.2},
  {16.9, 20.2, 20.6},
  {17, 19.1, 21.4},
  {18.2, 19.4, 21.9},
  {18.1, 20.5, 22.8},
  {17.2, 20, 22.2},
  {16, 19, 21.5},
  {15.1, 17.2, 20.1},
  {13.6, 15.8, 18.9},
  {12.6, 15.5, 16.8},
  {13.4, 14.6, 15.5},
  {13.8, 14.2, 14.4},
  {12.1, 13.5, 13.8},
  {10.7, 13, 13},
  {10.3, 12.3, 12},
  {10, 11.6, 11.5},
  {9.9, 11.2, 10.8},
  {11.6, 11.6, 10.7},
  {15.2, 12.2, 11.5},
  {16.4, 13.8, 14.6},
  {17.5, 16.4, 17.4},
  {18.2, 18.2, 20.3},
  {19.2, 20.3, 22.1},
  {20, 21.7, 23.8},
  {20.7, 22.3, 23.8},
  {21.1, 22.8, 23.7},
  {21.1, 23, 24},
  {20.6, 23.2, 24.1},
  {19.9, 22.4, 23.4},
  {19, 21.3, 22.7},
  {17.6, 20.6, 22.4},
  {17, 19, 21.4},
  {16.2, 17.6, 19.2},
  {16.3, 17.4, 17.3},
  {15.6, 17.5, 15.8},
  {14.8, 17, 14.7},
  {13.4, 15.8, 13.9},
  {11.9, 15.3, 13.2},
  {11.6, 15, 12.7},
  {11.5, 14.1, 12.4},
  {12.2, 13.7, 12},
  {13.2, 14.2, 12.2},
  {15.1, 15.1, 12.9},
  {17.6, 16.3, 14.7},
  {18, 17.1, 17.6},
  {18, 17.2, 18.9},
  {17.6, 17.9, 20.3},
  {20.1, 19.8, 22.5},
  {20.6, 21.5, 23.2},
  {19.7, 21.1, 23.1},
  {20.2, 21.4, 23.5},
  {20, 21.3, 23},
  {19.7, 21.1, 23.3},
  {19.5, 20.8, 23},
  {18.5, 20.9, 22.7},
  {17.4, 18.5, 21.5},
  {16.9, 17, 18.9},
  {15.4, 16.9, 17},
  {15, 16.9, 15.8},
  {14.3, 16.1, 15.1},
  {14.7, 15.6, 14.7},
  {14.7, 15.4, 14.5},
  {13.9, 14.2, 13.8},
  {14.5, 13.8, 13.3},
  {13.6, 13.9, 13.1},
  {13.5, 13.5, 13.5},
  {14.4, 13.9, 14.3},
  {15.3, 14.7, 16.2},
  {16.3, 16.9, 19.3},
  {17.3, 18.4, 21.4},
  {19, 20.2, 23.7},
  {19.9, 21.8, 23.7},
  {19.2, 21.5, 22.1},
  {17.8, 20.3, 21.1},
  {18.4, 20, 21.3},
  {17.7, 19.4, 21.4},
  {17.2, 19.1, 21.4},
  {16.2, 18, 21.3},
  {15.2, 17.4, 20.6},
  {14.6, 16.6, 20.1},
  {13.9, 16.2, 19.2},
  {13.4, 15.2, 18.5},
  {13.1, 14.1, 18.1},
  {13.2, 13.3, 17.9},
  {13.4, 13, 17.3},
  {13, 12.5, 15.6},
  {11.2, 12.9, 14.5},
  {10.1, 12.5, 13.9},
  {9.9, 12.1, 13.4},
  {10, 12.1, 13.1},
  {10.9, 12.8, 13.2},
  {11.8, 13.6, 13.7},
  {13.1, 14.6, 14.5},
  {15.2, 16.1, 16.1},
  {15.5, 17.4, 18.3},
  {16.3, 17.9, 20.3},
  {14.7, 17.9, 19.2},
  {14.8, 18, 20.1},
  {16.1, 17.6, 20},
  {16.4, 18.3, 20.3},
  {16.8, 18.6, 20.2},
  {15.9, 18.2, 19.1},
  {14, 16.6, 18.6},
  {13.5, 15.6, 17.6},
  {12.6, 14, 16.4},
  {11.8, 12.9, 15},
  {10.8, 12.8, 13.7},
  {10.5, 12.8, 12.7},
  {10.4, 12.1, 12},
  {10.6, 11.5, 11.6},
  {11.4, 11.8, 11.8},
  {11.2, 11.3, 11.7},
  {9.6, 11.6, 11.2},
  {10.7, 12, 11.2},
  {13, 12.5, 11.9},
  {13.1, 14, 12.3},
  {15, 16, 13.9},
  {16, 17.6, 17.1},
  {17.3, 18.7, 19.9},
  {18.2, 18.6, 21.4},
  {18.4, 19.6, 22.5},
  {16.6, 21.3, 22.1},
  {17.7, 20.9, 22.7},
  {18.4, 20.2, 23.5},
  {18, 19.7, 23.3},
  {16.8, 18.4, 22.7},
  {14.5, 16.3, 21.3},
  {13.3, 13.5, 19.4},
  {11.5, 11.9, 17.3},
  {10.3, 10.9, 15.7},
  {9.2, 10.3, 14.6},
  {7.9, 9.5, 13.7},
  {7.2, 9, 12.4},
  {7, 8.4, 11.3},
  {6.9, 8, 8.8},
  {6.3, 7.2, 7.9},
  {5.8, 6.7, 6.3},
  {5.9, 6.3, 5.5},
  {9, 7.3, 6.4},
  {9.6, 9.2, 10},
  {10.7, 11.5, 12.7},
  {11.7, 12.8, 15.8},
  {13.3, 14, 16.5},
  {14.8, 15.1, 17.5},
  {15.3, 16, 18.3},
  {15.5, 16.7, 19.1},
  {15.9, 16.9, 19.4},
  {15.5, 16.7, 19.4},
  {15.3, 16.3, 19.4},
  {14.6, 15.6, 18.8},
  {13.4, 14.5, 18.2},
  {12, 12.7, 17.1},
  {10.1, 11.9, 16},
  {9.7, 11.1, 15.3},
  {8.9, 9.6, 14.5},
  {8.7, 8.7, 12.1},
  {7.6, 8.2, 10.2},
  {6, 7.4, 8.5},
  {5.6, 8, 7.5},
  {5, 9, 6},
  {5.2, 8.9, 5.3},
  {7.1, 7.7, 5},
  {9.4, 7.6, 7},
  {10.4, 9.9, 10.2},
  {11.9, 11.9, 13.2},
  {12.4, 13.4, 15.7},
  {13.2, 14.3, 16.5},
  {14.2, 15.2, 17.9},
  {14.8, 15.9, 18.4},
  {14.9, 16.1, 19},
  {14.8, 16.3, 18.4},
  {14.1, 16.3, 17.8},
  {14.2, 15.8, 18},
  {13.2, 15.4, 17.7},
  {11.4, 14.1, 17.6},
  {10.9, 12, 16.5},
  {10.1, 10.7, 15.4},
  {9.7, 10.1, 15},
  {9.8, 9.6, 13.8},
  {9.2, 9.4, 11.6},
  {6.8, 8.9, 8.8},
  {4.6, 7.8, 7.1},
  {4.6, 7.7, 5.9},
  {4.6, 6.9, 4.8},
  {6.4, 6.1, 3.9},
  {7.5, 6.1, 3.6},
  {9.5, 6.8, 5.5},
  {9.8, 8.9, 8.6},
  {11, 11.8, 11.8},
  {12.5, 13.9, 15.6},
  {14, 15.4, 17.6},
  {15, 16.7, 18.7},
  {16, 18, 20.1},
  {16.7, 19, 21.1},
  {16.5, 19.2, 21.9},
  {16.4, 19.5, 21.3},
  {15.6, 19.5, 20.3},
  {15, 19.1, 19.9},
  {13.5, 17.9, 18.3},
  {12.4, 15.9, 15.4},
  {11.3, 13.6, 14.1},
  {9.2, 12.1, 13.2},
  {8.4, 12.1, 12.5},
  {8.9, 11.7, 11.2},
  {9.3, 10.1, 11},
  {9, 9.6, 10.9},
  {8.6, 8.8, 10.6},
  {7.8, 8.7, 9.8},
  {7.7, 8.3, 8.5},
  {8.1, 8.7, 7.7},
  {11.5, 9.6, 8.8},
  {12.4, 10.8, 12.2},
  {13.3, 12.4, 15.1},
  {14.8, 13.8, 16.6},
  {15.7, 16.3, 18.8},
  {15.2, 17.8, 19.2},
  {15.7, 18.4, 19.5},
  {15, 18.5, 20.5},
  {14.8, 17.9, 20.5},
  {15.5, 18.1, 20.5},
  {15.4, 18.4, 20.2},
  {15.1, 18.1, 19.6},
  {14.7, 17.1, 19.2},
  {14, 16.3, 18.7},
  {13.1, 15.5, 17.9},
  {13.2, 15, 16.5},
  {13.2, 15.3, 15.4},
  {12.5, 14.9, 16.3},
  {11.9, 14.2, 15.7},
  {11.6, 13.7, 14.5},
  {11.3, 13.7, 13.8},
  {10.7, 12.9, 12.5},
  {10.2, 12.1, 11.4},
  {10.5, 12.9, 11},
  {11.3, 13.2, 11.5},
  {11.3, 13.7, 14},
  {13, 14.4, 15.7},
  {15.4, 15.3, 17.6},
  {15.2, 16.4, 18.8},
  {14.8, 17.7, 19.3},
  {14.8, 17.8, 17.8},
  {13.3, 16.7, 16},
  {14.2, 16.1, 17},
  {15.3, 17.1, 17.8},
  {15.9, 17.7, 19},
  {15.7, 18.2, 19.9},
  {15.1, 17.4, 19},
  {14.8, 16.1, 16.9},
  {14.5, 15.5, 15},
  {14.4, 15.3, 13.9},
  {14, 15.1, 13.4},
  {13.4, 14.7, 13.4},
  {12.7, 14.4, 13.1},
  {11.8, 14.1, 12.5},
  {11.5, 14.1, 12.1},
  {11.6, 13.8, 11.8},
  {11.5, 13.7, 12.1},
  {11.8, 13.7, 12.4},
  {12.1, 13.8, 13},
  {12.3, 14, 13.6},
  {13.5, 14.9, 14.9},
  {15.4, 16.5, 16.8},
  {16.3, 16.6, 17.7},
  {17.2, 18.1, 19.7},
  {17.9, 20.1, 20.7},
  {18.2, 20.4, 19.8},
  {18, 19.8, 20.3},
  {17.3, 20.1, 20.4},
  {16.8, 20, 20.1},
  {16.1, 19.1, 20},
  {15.7, 18, 19.7},
  {15.3, 17.5, 18.9},
  {14.1, 16.3, 17},
  {14.6, 15.5, 15.9},
  {12.7, 15.5, 14.6},
  {12.2, 15.8, 14.1},
  {11.8, 15.2, 13.4},
  {11.6, 15.2, 12.9},
  {12.7, 15, 12.8},
  {12.7, 14.3, 12.9},
  {13.5, 13.5, 13.1},
  {14, 14.2, 13.4},
  {14.7, 14.9, 13.8},
  {13.9, 14.7, 14.3},
  {13.2, 14.2, 14.6},
  {13.3, 14.3, 14.3},
  {13.3, 13.9, 14.4},
  {13.3, 14.8, 14.6},
  {13.3, 14.5, 14.8},
  {13.7, 14.4, 15.1},
  {13.3, 14.3, 15.2},
  {13.4, 14.6, 15.4},
  {13, 14.5, 15.5},
  {12.9, 14.3, 15.5},
  {12.6, 13.7, 15.5},
  {12.6, 13.5, 14.8},
  {12.4, 13.4, 14.5},
  {12.4, 13.2, 14.5},
  {12.3, 13.2, 14.4},
  {12.3, 13.1, 14.4},
  {12.3, 13.1, 14.3},
  {11.7, 13, 14.1},
  {11.7, 13, 14},
  {10.5, 12.9, 14},
  {10.7, 12.9, 13.8},
  {11.3, 13.1, 13.9},
  {13, 13.5, 14.2},
  {14.6, 14.3, 14.2},
  {15.6, 16, 15.4},
  {16.2, 17.1, 18.8},
  {17.2, 17.3, 19.9},
  {17.5, 19, 21.9},
  {17.7, 20, 22.2},
  {17.9, 20, 21},
  {16.3, 20.6, 21.8},
  {16.7, _, 19.9},
  {16.9, _, 20.3},
  {17.1, _, 19},
  {15.9, _, 18.9},
  {14.4, _, 18.2},
  {13.8, _, 17.1},
  {13.4, _, 15.9},
  {13.8, _, 15.2},
  {14.2, _, 15.2},
  {14.1, _, 15},
  {13.4, _, 14.8},
  {12.8, _, 14.6},
  {13.3, _, 14.3},
  {13.5, _, 13.8},
  {13.7, _, 14.1},
  {14.7, _, 14.5},
  {15.7, _, 15},
  {17.9, _, 16.6},
  {18.8, _, 19.5},
  {20.1, _, 22.8},
  {20.9, _, 25.1},
  {22.4, _, 26.7},
  {22.8, _, 27.8},
  {23, _, 26.8},
  {22.7, _, 26.1},
  {22.5, _, 25.6},
  {21.7, _, 25.3},
  {19.6, _, 24.8},
  {17.7, _, 23.3},
  {16.6, _, 20.4},
  {15.7, _, 18.4},
  {15.5, _, 17.1},
  {15.6, _, 16.3},
  {15.4, _, 15.6},
  {14.6, _, 14.8},
  {14.4, _, 14.3},
  {13.8, _, 13.8},
  {13.6, _, 13.4},
  {14.6, _, 13.3},
  {17.6, _, 14.3},
  {18.7, _, 16.6},
  {18.9, _, 20.1},
  {20.1, _, 22.2},
  {21.4, _, 24.4},
  {22.7, _, 26.3},
  {23.2, _, 27.5},
  {22.6, _, 25.7},
  {22.6, _, 25.3},
  {22.9, _, 26.3},
  {21.8, _, 25.8},
  {20.8, _, 24.9},
  {19.6, _, 23.9},
  {18.8, _, 22.5},
  {16.5, _, 20.6},
  {16.1, _, 18.7},
  {15.6, _, 17.6},
  {15.5, _, 16.8},
  {16.1, _, 16.3},
  {15.8, _, 15.8},
  {16.1, _, 15},
  {15.4, _, 14.2},
  {14.6, _, 13.7},
  {16.4, _, 13.4},
  {19.1, _, 14.5},
  {20.1, _, 17.9},
  {21, _, 19.3},
  {22.8, _, 21.9},
  {24, _, 24.9},
  {24.6, _, 27.2},
  {25.5, _, 29.4},
  {26, _, 30},
  {25.6, _, 29.8},
  {24.8, _, 28.8},
  {24.6, _, 28.4},
  {24, _, 27.9},
  {22.5, _, 27.3},
  {21.1, _, 25.9},
  {19.3, _, 22.9},
  {19, _, 21},
  {19.1, _, 19.9},
  {18.2, _, 19.2},
  {18.4, _, 18.2},
  {18.4, _, 17.9},
  {18.4, _, 17.6},
  {18.3, _, 17.5},
  {18.1, _, 17.6},
  {18, _, 17.9},
  {18.8, _, 18.7},
  {19.6, _, 19.7},
  {20.3, _, 21.7},
  {21, _, 24},
  {21.8, _, 25.9},
  {22.2, _, 25.7},
  {22.6, _, 25.7},
  {22.7, _, 26.2},
  {22.9, _, 26.7},
  {23.5, _, 26.7},
  {22.8, _, 27.2},
  {21.1, _, 26},
  {20, _, 24.8},
  {19.1, _, 23.8},
  {18.8, _, 22.4},
  {17.8, _, 19.7},
  {17.6, _, 18.6},
  {16.5, _, 17.8},
  {16, _, 17.3},
  {14.5, _, 17},
  {14, _, 16.6},
  {14.2, _, 16.3},
  {14.2, _, 15.8},
  {14.9, _, 15.5},
  {17.5, _, 16.9},
  {18.2, _, 19.1},
  {19.4, _, 21.5},
  {20.3, _, 23.5},
  {21.7, _, 24.4},
  {22.3, _, 25.1},
  {22.6, _, 25.3},
  {22.9, _, 26},
  {22.6, _, 26.3},
  {22.4, _, 26.2},
  {22.1, _, 26.2},
  {21.3, _, 25.4},
  {20, _, 24.5},
  {19.6, _, 23.4},
  {19.4, _, 21.8},
  {19.2, _, 21},
  {18.6, _, 20.6},
  {17.5, _, 19.3},
  {17.3, _, 18},
  {17.4, _, 18.6},
  {15.9, _, 18.1},
  {14.1, _, 17.5},
  {13.7, _, 17.2},
  {15.2, _, 16.6},
  {17.5, _, 17.8},
  {19, _, 20.1},
  {20.5, _, 22.9},
  {21.4, _, 24.2},
  {22.7, _, 25.9},
  {23.7, _, 27.7},
  {24.3, _, 28.2},
  {24.9, _, 27.5},
  {24.7, 27.4, 27.2},
  {23.2, 26.8, 28.4},
  {23.4, 25.9, 28.1},
  {23, 25.3, 26.4},
  {21.2, 24.1, 24.9},
  {20.1, 23, 24},
  {19.8, 21.4, 21.8},
  {19.4, 20.5, 20.3},
  {17.9, 19.9, 19.1},
  {17.9, 19.6, 18.5},
  {16.7, 18.9, 18},
  {16, 18.6, 17.2},
  {15.8, 17.6, 16.7},
  {15.8, 17.2, 16.2},
  {15.3, 17.2, 15.4},
  {15.9, 17.2, 14.9},
  {19.8, 17.4, 15.8},
  {21.2, 19.7, 19.3},
  {21.7, 22.9, 21.9},
  {22.3, 25, 24.3},
  {24.6, 25.9, 27.4},
  {25.7, 26.9, 29.7},
  {26.2, 28.9, 29.3},
  {26.5, 29.7, 28.9},
  {25.8, 28.6, 29.9},
  {25.6, 28.1, 29.7},
  {25.1, 27, 30},
  {24.3, 26.4, 29},
  {23.2, 25.4, 27.8},
  {21.8, 24.1, 26.1},
  {19.6, 23.1, 23.5},
  {19.2, 22.7, 21.4},
  {20.3, 22.5, 20.2},
  {20.5, 21.7, 19.1},
  {19.6, 21, 18.4},
  {18, 20.3, 17.6},
  {16.6, 19.6, 17.1},
  {16, 18.8, 16.5},
  {16.2, 18.2, 16},
  {17.4, 18.4, 16},
  {20.4, 18.9, 17.1},
  {22, 19.9, 20.1},
  {22.7, 22.9, 22.7},
  {23.9, 24.7, 25.1},
  {25.1, 25.4, 27.5},
  {26.2, 27, 29.4},
  {26.4, 29.2, 30},
  {27.3, 30.3, 29.9},
  {26.3, 29.9, 29.5},
  {24.1, 28.5, 28.9},
  {23, 26.4, 26.9},
  {23.3, 26.3, 25.1},
  {23.3, 25.8, 25.6},
  {22.8, 24.5, 24.4},
  {22.3, 23.7, 23},
  {22, 23.7, 21.6},
  {21.9, 23.7, 20.7},
  {21.2, 23.5, 20.2},
  {20.9, 23, 19.9},
  {20.9, 22.5, 19.6},
  {20.1, 21.4, 19.5},
  {19.5, 21.1, 19.1},
  {19.8, 21.9, 19},
  {19.9, 21.7, 19.3},
  {20.5, 21.9, 19.8},
  {21.6, 22.8, 20.9},
  {22.5, 23.6, 22.5},
  {23.7, 24.8, 24.6},
  {24.6, 26.1, 27.4},
  {25.2, 27.3, 28.2},
  {25.2, 27.7, 27.9},
  {25.4, 26.4, 27.9},
  {25.8, 25.6, 27.5},
  {25.5, 24.9, 26.3},
  {22.9, 24, 23},
  {22.4, 23, 21.2},
  {21.7, 21, 20.2},
  {20.1, 18.9, 20},
  {18.9, 18.6, 19.4},
  {18.4, 19.6, 18.7},
  {18.3, 18.7, 18.2},
  {17.6, 18.6, 17.8},
  {16.8, 17.5, 17.4},
  {16.1, 17, 17},
  {15.8, 16.7, 16.8},
  {15.4, 16.4, 16.9},
  {15.5, 16, 17.1},
  {16.2, 16.2, 17.3},
  {17.7, 16.9, 17.4},
  {18.7, 18, 17.8},
  {20.3, 19.5, 18.7},
  {21.6, 21.1, 20.8},
  {23.4, 23.1, 23.5},
  {24.4, 25.4, 26.3},
  {25.6, 27.1, 28.2},
  {26.3, 27.9, 28.6},
  {25.5, 27.6, 28.2},
  {25.6, 25.3, 26.8},
  {24, 24.4, 23.4},
  {21.8, 19.7, 20.1},
  {21.7, 18.1, 18.6},
  {21.4, 17.6, 18.5},
  {19.9, 17.2, 18.3},
  {18.5, 17.5, 17.7},
  {17.6, 17.4, 17.2},
  {17.1, 17.1, 16.8},
  {17.1, 16.6, 16.6},
  {16.9, 16.8, 16.7},
  {15.9, 16.4, 16.7},
  {15.8, 16.4, 16.3},
  {15.3, 16.3, 16.2},
  {15.9, 16.1, 16},
  {19.6, 16.4, 16.1},
  {20.8, 17.6, 16.8},
  {21.9, 21.4, 19.4},
  {23.5, 23.5, 21.9},
  {24.9, 25.8, 24.7},
  {26, 28.3, 27.6},
  {27.4, 29.8, 29.7},
  {28.1, 30.8, 30.7},
  {27.2, 31.5, 30.3},
  {27, 30.6, 30.2},
  {26.2, 29.3, 29.9},
  {25.1, 28.1, 29.3},
  {23.8, 27.3, 28.3},
  {23, 25.6, 26.6},
  {22.7, 24, 23.3},
  {22, 23.5, 21.2},
  {21.4, 22.9, 19.9},
  {20.2, 21.8, 19},
  {20.1, 21, 18.2},
  {19.9, 20.9, 17.7},
  {18.3, 20.3, 17.3},
  {17.4, 19.7, 16.8},
  {17.1, 18.8, 16.4},
  {18, 19.2, 16.3},
  {20.6, 19.9, 17.3},
  {21.7, 20.7, 19.7},
  {23, 22.3, 22.3},
  {24, 24, 24.8},
  {25.3, 26, 27.2},
  {26.6, 27.8, 29},
  {26.9, 29.4, 29.9},
  {27.4, 29.9, 29.6},
  {25.2, 29.7, 29.7},
  {22.6, 29, 28.4},
  {21.3, 28.1, 27.9},
  {21.5, 27.6, 27.9},
  {20.9, 26.6, 27.7},
  {19.7, 25.2, 26.1},
  {19.7, 23.5, 23.5},
  {19.5, 22.5, 22},
  {19.6, 22.5, 21.1},
  {20, 22.1, 20.5},
  {19.7, 21.1, 19.8},
  {19.6, 20.2, 19.3},
  {19.5, 20.2, 19.1},
  {19.4, 20, 19.1},
  {19.4, 19.6, 18.8},
  {19.7, 19.4, 19.1},
  {21.1, 20, 20.4},
  {22, 21, 22.5},
  {22.9, 23.9, 24.7},
  {24.5, 25.5, 26.1},
  {25.6, 26.8, 28.2},
  {26.8, 28.1, 29.9},
  {27.4, 29.7, 31.5},
  {28.1, 30.9, 32.5},
  {25.2, 30.2, 30.1},
  {24.1, 29.5, 29.2},
  {24.2, 28.7, 29.3},
  {24.5, 28.2, 28.8},
  {24, 27.4, 27.4},
  {22.4, 25.9, 26.1},
  {22.1, 24.6, 23.7},
  {21.4, 24.3, 22.1},
  {22, 23.8, 21.4},
  {20.2, 22.5, 20.2},
  {19.9, 22.1, 19.8},
  {19, 22.5, 19.2},
  {19.3, 21.8, 18.7},
  {19.3, 21.2, 18.3},
  {19.9, 21, 18.3},
  {20.3, 21.3, 18.8},
  {21.7, 21.7, 19.4},
  {23.2, 22.4, 20.9},
  {23.4, 23.3, 23.7},
  {24.9, 24.2, 25.8},
  {24, 25.2, 26.7},
  {19.7, 23.2, 23.7},
  {18.9, 24.3, 21.8},
  {20.9, 26.2, 21.2},
  {20.5, 22.3, 21.4},
  {21.8, 20.6, 20.5},
  {23, 20.9, 21.3},
  {21.5, 19.3, 21.2},
  {18.9, 16.8, 20.7},
  {15.1, 16.7, 17.3},
  {15.1, 17, 16.9},
  {15.3, 16.6, 17.1},
  {15.2, 16.6, 17.2},
  {14.9, 16.4, 17.1},
  {14.8, 16.2, 17},
  {14.4, 15.8, 16.9},
  {13.8, 15.7, 16.4},
  {13, 15.9, 16.4},
  {12.8, 16, 15.7},
  {13.8, 16, 15.7},
  {15.9, 16.1, 16.3},
  {17.1, 16.7, 17},
  {18.3, 18.2, 19.1},
  {19.3, 19.4, 21.2},
  {20.8, 20.9, 22.9},
  {22.2, 22.7, 25},
  {23.5, 24.4, 27.3},
  {24.7, 26.3, 27.2},
  {24.4, 26.5, 25.6},
  {23.2, 25.8, 24.8},
  {22.8, 25.4, 22.3},
  {23, 24.6, 23.4},
  {21.3, 23.7, 24.8},
  {20.3, 21.8, 22.7},
  {17.8, 21.3, 20.1},
  {18.6, 20.9, 18.5},
  {18.7, 20.3, 17.8},
  {18.4, 19.7, 17.4},
  {17.6, 19.8, 17.5},
  {18, 19, 17.2},
  {18.1, 17.5, 17.1},
  {16.9, 16.7, 17.1},
  {16.7, 15.3, 17.1},
  {15.3, 14.8, 17.1},
  {14.3, 14.8, 17.2},
  {14.4, 15, 17.2},
  {14.3, 15.6, 17.6},
  {14.5, 14.9, 17.9},
  {14.5, 14, 17.5},
  {14.9, 14.2, 18.3},
  {15.7, 15.8, 19.2},
  {17, 17, 21.5},
  {18.2, 19.3, 22.7},
  {19.2, 21, 23.7},
  {19.9, 21.6, 24.4},
  {19.3, 21, 22.9},
  {17.1, 19.9, 21.7},
  {15.4, 17.8, 19.8},
  {14.1, 17.3, 17},
  {12.8, 16.3, 15.3},
  {13.3, 15.5, 14.1},
  {13.5, 14.9, 13.4},
  {13.4, 14.1, 13.1},
  {12.9, 14, 12.6},
  {11.9, 14.6, 11.7},
  {12.2, 14.7, 11.1},
  {12.2, 14.5, 10.6},
  {13.9, 14.3, 10.3},
  {16.3, 14.5, 11},
  {16.8, 15.2, 14},
  {17.2, 17.9, 17.7},
  {18.4, 19.6, 21.4},
  {19.9, 21.7, 23.6},
  {21.4, 23, 24.8},
  {22.4, 24, 25.4},
  {22.8, 24.7, 25.8},
  {23.3, 25.5, 26.7},
  {24, 26.1, 27.1},
  {23.7, 25.9, 27.5},
  {22.5, 25.3, 26.6},
  {19.5, 24.5, 24.9},
  {17.4, 22.2, 22.7},
  {16, 19.9, 18},
  {15.7, 18.7, 16.3},
  {16.9, 17.8, 14.9},
  {16, 17.4, 14.1},
  {14.8, 16.7, 13.2},
  {14.2, 16.3, 12.5},
  {13.9, 15.7, 11.8},
  {13, 14.9, 11.3},
  {12.1, 14.6, 10.7},
  {13.8, 14.3, 10.4},
  {17.7, 14.9, 11.4},
  {18, 15.9, 14.9},
  {18.8, 18.9, 18.4},
  {19.6, 21.3, 20.8},
  {20.6, 21.5, 23.8},
  {21.4, 23, 25.3},
  {22.1, 24.8, 25.7},
  {22.1, 25.5, 25.8},
  {22, 25.6, 25.9},
  {22, 25.4, 25.8},
  {21.9, 25, 25.6},
  {21.4, 24.2, 25.2},
  {19.9, 23.3, 24.3},
  {19, 21.6, 22.9},
  {18.2, 20.7, 20.6},
  {18.7, 19.9, 19.3},
  {17.8, 19.8, 18.4},
  {18, 19.3, 18.4},
  {17.6, 19.3, 18.3},
  {17, 19.6, 18.3},
  {16.9, 19.2, 18.2},
  {16.6, 19.1, 18},
  {15.9, 18.2, 17.9},
  {15.7, 17.8, 17.7},
  {18, 17.5, 18.1},
  {18.9, 18.7, 19.3},
  {19.9, 21.2, 22.1},
  {21, 22.1, 23.3},
  {21.2, 23.1, 23.8},
  {21.6, 24.1, 24.8},
  {21.5, 24.8, 25.4},
  {21.9, 25.1, 25.8},
  {21.9, 25.2, 25.6},
  {20.9, 25.2, 25.2},
  {21.1, 24.3, 24.9},
  {21, 23.8, 24.9},
  {20.2, 22.7, 24},
  {18.4, 21.3, 23.4},
  {19.3, 19.4, 21.9},
  {19.1, 19.7, 19.9},
  {19.1, 19.9, 19.6},
  {18.5, 19.6, 19.3},
  {17.3, 18, 19},
  {15.2, 16.7, 17.7},
  {14.1, 16.5, 17.4},
  {13.3, 15.8, 17.2},
  {13.6, 14.9, 17},
  {13.9, 14.9, 16.7},
  {14.5, 14.8, 16.7},
  {14.3, 15.1, 17},
  {13.8, 13.5, 17},
  {14.2, 11.5, 17},
  {12.7, 10.9, 15.7},
  {10.5, 10.7, 14.4},
  {10.7, 11, 13.8},
  {11.3, 13, 16.2},
  {13, 15.3, 18.3},
  {15.2, 16.1, 19.4},
  {16.3, 17.1, 19.5},
  {15.8, 17.6, 20.1},
  {13.4, 17.3, 19},
  {11.5, 15.5, 16.5},
  {10.7, 13.4, 14.2},
  {10.7, 12.8, 12.7},
  {10.6, 11.9, 11.5},
  {9.9, 11.2, 10.6},
  {8.9, 11.1, 9.8},
  {8.5, 10.5, 9.2},
  {7.7, 9.9, 8.5},
  {7.4, 9.2, 8},
  {7.1, 9.1, 7.5},
  {8.4, 9.3, 7.2},
  {12.4, 9.5, 7.9},
  {13.7, 11.2, 10.4},
  {14, 14.1, 14.1},
  {14.9, 15.2, 16.9},
  {15.9, 16.3, 19.8},
  {17.2, 18.8, 21.2},
  {17.9, 20, 21.2},
  {18.5, 20.7, 21.7},
  {18.8, 21.3, 21.8},
  {18.9, 21.1, 21.9},
  {18.2, 20.4, 21.4},
  {17.4, 19.8, 21.1},
  {16.4, 18.6, 20.6},
  {15.4, 17.5, 18.7},
  {15.4, 16.3, 17.6},
  {15.2, 15.7, 15.7},
  {13.8, 16, 14.3},
  {12.2, 15.5, 13.2},
  {11.6, 14.6, 12.3},
  {11.5, 14, 11.6},
  {12.6, 13.9, 11.2},
  {12.6, 13.7, 11.9},
  {12.3, 13.4, 12},
  {12.8, 13.3, 12},
  {13.7, 13.8, 12.9},
  {14.3, 15.1, 14.5},
  {15.1, 15.8, 15.6},
  {15.7, 16.2, 17.5},
  {14.8, 16.7, 17.7},
  {13.9, 16.2, 16},
  {14.1, 15, 15},
  {14.9, 14.6, 15.3},
  {15, 14.6, 16.3},
  {16.2, 15.7, 17.1},
  {15.1, 15.8, 17.3},
  {14.5, 15.1, 17.1},
  {13.8, 14.2, 17.2},
  {12.7, 13.9, 16.7},
  {12, 13.6, 16.3},
  {12.1, 13.2, 15.6},
  {12, 10.6, 15},
  {11.6, 9.9, 13.9},
  {10.1, 9.6, 12.9},
  {9.2, 9.4, 12.3},
  {8.7, 9.3, 12},
  {8.4, 9.2, 11.7},
  {8.1, 9.1, 11.4},
  {8.4, 9.1, 11.5},
  {9.5, 9.3, 11.8},
  {11.5, 10.2, 12.8},
  {12.6, 12.1, 15.1},
  {13.9, 14, 17.1},
  {15.5, 17, 19.2},
  {17.1, 18.8, 21},
  {18.3, 20.2, 22},
  {19.1, 21.5, 22},
  {19.3, 20.5, 21.3},
  {18.7, 19.7, 19.4},
  {15.5, 20.3, 19.3},
  {14.6, 19.2, 18.4},
  {13.6, 18.3, 17.9},
  {13.1, 16.9, 17.5},
  {11.9, 15, 15.5},
  {12.1, 14.5, 13.7},
  {12.6, 13.8, 12.4},
  {11.9, 12.7, 11.6},
  {12.4, 13.2, 11.1},
  {12.4, 13.3, 11.5},
  {12.1, 13.2, 11.8},
  {12, 12.7, 11.6},
  {12.1, 11.9, 11.2},
  {12.3, 11.8, 11.4},
  {12.6, 12.2, 11.9},
  {12.6, 12.4, 12.4},
  {12.8, 13.3, 13},
  {13.5, 14.1, 13.6},
  {13.9, 14.3, 15.1},
  {14.9, 15, 16.6},
  {15.2, 16.3, 18.3},
  {15.7, 16.8, 19.6},
  {15.8, 17.3, 20.3},
  {16.5, 18, 21},
  {16.3, 18.3, 20.3},
  {15.9, 16.7, 20.5},
  {15.1, 15.2, 19.1},
  {14.5, 14.3, 18.5},
  {13.6, 13.4, 17.1},
  {12.8, 13.1, 15.9},
  {11.6, 13.3, 15},
  {11.6, 13.5, 14},
  {11.2, 13, 14},
  {11, 12.8, 13.7},
  {10, 12.8, 12.8},
  {10.5, 12.4, 12.5},
  {10.9, 12.4, 12},
  {11.9, 12.7, 11.8},
  {12.6, 12.6, 12.6},
  {13.8, 13.7, 15.4},
  {15.4, 16.4, 17.4},
  {16, 18.2, 19.9},
  {16.8, 19.5, 21.5},
  {17.4, 19.1, 22.4},
  {18.4, 19.2, 22.3},
  {18, 18.1, 23},
  {16.9, 15.5, 22.1},
  {16.1, 14.4, 21.4},
  {15.1, 15, 19},
  {15.6, 16.5, 18.1},
  {14.7, 15.8, 17.7},
  {13.8, 14.3, 16.7},
  {13.1, 13.8, 15.9},
  {12.9, 13.2, 15.1},
  {12.6, 13.2, 14.7},
  {12, 13.1, 14.5},
  {11.9, 13.1, 14.2},
  {11.7, 13.1, 14},
  {11.4, 12.8, 13.9},
  {11.2, 12.6, 13.7},
  {11.3, 12.4, 13.5},
  {11.4, 12.5, 13.3},
  {12.6, 12.7, 13.6},
  {14.4, 13.3, 14.4},
  {16.5, 15.4, 16.8},
  {16.8, 15.5, 19.5},
  {17.2, 16.5, 20.9},
  {18.7, 19.1, 22.7},
  {20.1, 21.2, 24.2},
  {19.8, 22.4, 25.5},
  {20.7, 22.6, 25.4},
  {20.5, 22, 25.8},
  {19.4, 21.2, 25},
  {18.8, 20.8, 23.3},
  {18.2, 20.1, 22.6},
  {16.7, 19, 21.4},
  {15.5, 18.4, 19.1},
  {14.3, 17.5, 17},
  {14.7, 17.2, 15.4},
  {14.3, 16.7, 14.1},
  {15, 15.3, 13.4},
  {15, 15.1, 12.4},
  {14.6, 15.2, 12.1},
  {13.6, 14.3, 11.8},
  {13.9, 14, 11},
  {14, 14.2, 10.5},
  {16.5, 14.9, 11.5},
  {16.8, 16.6, 13.3},
  {18.4, 18.9, 16.1},
  {18.3, 20.7, 18.1},
  {20.7, _, 21.7},
  {22, 22.3, 23.9},
  {21.6, 22.7, 25.6},
  {22.3, 23.9, 25.8},
  {22.5, 24.6, 27.6},
  {22.4, 24.8, 25.8},
  {20.1, 23.4, 22.4},
  {19.3, 22.6, 21.4},
  {18.6, 21, 21.2},
  {16.7, 19.5, 20.1},
  {15.2, 18.3, 17.9},
  {15.1, 17, 16.1},
  {15.2, 16.6, 15},
  {14.5, 17, 13.8},
  {14, 17.1, 13},
  {13.6, 16.4, 12.5},
  {13.3, 15.8, 12.2},
  {12.6, 15.2, 11.6},
  {12.8, 14.4, 11.1},
  {13.2, 14.7, 11},
  {14.4, 15, 12},
  {17.1, 15.9, 14.2},
  {18.7, 18.6, 17.1},
  {19, 20, 20.2},
  {20.3, 21.9, 22.1},
  {21.1, 23.4, 23.8},
  {21.8, 24.7, 26.2},
  {22.4, 26.2, 26},
  {22.4, 26.2, 26},
  {21.9, 26.1, 25.8},
  {21.7, 25.2, 25.3},
  {20.9, 24.1, 24.8},
  {19.7, 22.9, 24},
  {19.1, 21.3, 22.5},
  {18.7, 19.7, 21.3},
  {18, 19.4, 19.1},
  {17.7, 18.8, 17.3},
  {16.2, 17.5, 16.2},
  {14.8, 17.2, 15.2},
  {14.3, 16.2, 14.5},
  {14.1, 15.3, 13.7},
  {14, 15.4, 13.2},
  {14.1, 15.2, 12.6},
  {14.2, 14.8, 12.4},
  {17.4, 15, 13.3},
  {18.2, 16.1, 15.7},
  {18.8, 19.1, 19.5},
  {19.9, 21.5, 21.7},
  {21.4, 23.3, 24.2},
  {22.6, 24.1, 26.3},
  {23.6, 25.5, 27.8},
  {24.2, 26.8, 28.4},
  {24.1, 28, 28},
  {23.5, 27.7, 27.3},
  {23.4, 26.6, 27},
  {22.4, 25.6, 26.5},
  {21.1, 24.6, 25.3},
  {20, 22.8, 23.8},
  {19.3, 21.6, 21.3},
  {18.7, 20.9, 18.7},
  {17.7, 19.9, 17.4},
  {16.5, 19, 16.5},
  {15.6, 18.3, 16.1},
  {15.7, 17.5, 15.6},
  {15.5, 17.3, 15},
  {15.5, 17, 14.6},
  {15, 16.7, 14.2},
  {15.9, 17.5, 14.7},
  {18.4, 18.4, 15.8},
  {20.3, 18.8, 18},
  {21.3, 20.1, 21.2},
  {22.3, 21.8, 23.3},
  {23.2, 23.6, 25.3},
  {23.8, 25.3, 27.1},
  {23.8, 26.4, 27.5},
  {24, 27.1, 27.7},
  {24, 27.4, 27.8},
  {24.1, 26.8, 27.8},
  {23.8, 26.4, 27.4},
  {22.9, 25.2, 26.1},
  {21.9, 24.3, 26.2},
  {20.5, 23.1, 23.3},
  {17.5, 21.4, 20.1},
  {17.9, 20.6, 18.7},
  {16.7, 20.5, 17.4},
  {16.2, 19.4, 16.6},
  {16.1, 18.1, 16},
  {16, 17.4, 15.4},
  {15.5, 17, 15.8},
  {15.5, 16.8, 15.8},
  {15.8, 16.6, 16.2},
  {16, 16.8, 16.4},
  {19.1, 17.1, 16.5},
  {19.9, 18.3, 16.8},
  {20.2, 20.4, 18.3},
  {20.3, 20.9, 19.6},
  {20.9, 21.1, 22.2},
  {23, 22.1, 23.3},
  {23.5, 23.4, 25.3},
  {25, 25.2, 27.7},
  {25.1, 26, 27.6},
  {25.1, 25, 28},
  {22.1, 23.8, 26.6},
  {21.5, 23.7, 24.7},
  {21, 23.2, 24},
  {19.3, 21.1, 21.8},
  {18.7, 20.3, 19.7},
  {18.2, 20, 18.5},
  {17.9, 18.7, 17.8},
  {18, 18.1, 17.5},
  {18.1, 17.5, 17.2},
  {18.1, 17.3, 16.3},
  {18.2, 17, 16.3},
  {17, 17.1, 16.3},
  {17.3, 16.8, 15.5},
  {16.7, 16.6, 15.2},
  {18.5, 17, 15.9},
  {19.9, 17.7, 17.2},
  {20.7, 19.7, 19.4},
  {21.4, 22.6, 22.8},
  {23.2, 24, 25.4},
  {23.9, 24.8, 27.2},
  {25, 26.6, 29},
  {25.9, 28.1, 28.5},
  {26.6, 29, 28},
  {26.4, 28.4, 28.2},
  {25.5, 27.4, 28.2},
  {24.1, 26.6, 28.3},
  {22.4, 25.4, 27.6},
  {21.5, 24.1, 25.7},
  {20.9, 23, 22.5},
  {20.4, 22.2, 20.9},
  {19.7, 22.2, 19.8},
  {19.4, 21.2, 18.9},
  {18.2, 21.4, 18.1},
  {17.3, 20.4, 17.6},
  {17.1, 19.4, 16.9},
  {17, 18.8, 16.6},
  {17.9, 19.7, 17.1},
  {18.2, 19.8, 17.7},
  {19.6, 20.2, 18.5},
  {21.2, 20.7, 19.7},
  {21.2, 22.1, 22.2},
  {21.9, 22.9, 24},
  {23.3, 24.6, 26.2},
  {24.4, 26.2, 27.7},
  {24.7, _, 27.3},
  {22.2, 25.5, 26.7},
  {22, 21, 24.4},
  {23, 21.6, 26.3},
  {23.4, 22.8, 26.5},
  {22.8, 22.3, 26.2},
  {22.2, 20.9, 25.5},
  {21.3, 20.9, 24.5},
  {19.7, 20.3, 22.5},
  {20.5, 19.4, 20.8},
  {20.7, 19.7, 20.5},
  {20.4, 18.2, 21.1},
  {19.3, 14.6, 20.6},
  {18.2, 13.1, 18.2},
  {12.7, 12.6, 16.2},
  {11.8, 12.5, 14.7},
  {11.1, 12.6, 13.9},
  {10.7, 12.6, 13.5},
  {11.9, 12.8, 13.8},
  {13.4, 13.9, 14.8},
  {15.7, 15.7, 17.7},
  {16.3, 17.7, 20},
  {18.1, 19.9, 21.6},
  {20.2, 21.4, 23.6},
  {21.8, 23.2, 25.4},
  {23.1, 24.3, 26.8},
  {24, 24.5, 27.9},
  {23.4, 22.2, 29},
  {21.5, 22.1, 26.5},
  {20.8, 23.8, 25},
  {19.2, 23.4, 24.5},
  {17.5, 20.1, 21.2},
  {16, 18.6, 19},
  {15.9, 17.5, 17},
  {15.8, 18.1, 15.7},
  {15.7, 17.9, 14.8},
  {15.7, 17.3, 14.4},
  {15.8, 16.5, 14},
  {15, 15.9, 14},
  {13.7, 15.5, 13.6},
  {13, 15, 12.8},
  {13.9, 14.3, 12.3},
  {17.5, 14.4, 12.7},
  {18.7, 15.3, 16.1},
  {19.1, 18.4, 18.7},
  {19.6, 21.1, 21.4},
  {21.1, 21.3, 24},
  {22.1, 23.1, 26},
  {22.9, 25, 26.5},
  {22.9, 25.8, 26.7},
  {22.7, 26.1, 26.3},
  {22.9, 25.9, 26.6},
  {22.5, 25.6, 26.4},
  {22, 24.4, 25.3},
  {20.9, 23.5, 24.4},
  {20.1, 22, 23},
  {18.8, 20.8, 19.7},
  {17.2, 20.6, 18.4},
  {16.4, 19.8, 17.2},
  {16.3, 18.7, 16.2},
  {16.8, 18.1, 15.5},
  {15.8, 17, 14.9},
  {15.3, 16.5, 14.6},
  {15.1, 15.9, 13.9},
  {14.3, 16.1, 13.3},
  {15, 16, 12.8},
  {18.1, 16.2, 13.7},
  {19.5, 16.7, 16.1},
  {19.4, 19.7, 19.3},
  {19.9, 21.6, 22.1},
  {21.6, 23, 24.9},
  {22.9, 24.2, 27.1},
  {23.9, 25.4, 28.1},
  {23.6, 26.3, 28.6},
  {20.7, 27.3, 26.6},
  {20.1, 27.1, 25.4},
  {20.9, 25.4, 26.1},
  {21.6, 24.4, 25.8},
  {20.1, 22.9, 25},
  {18.2, 21.5, 22.8},
  {16.6, 21, 19.8},
  {17.2, 20.2, 18.3},
  {18.2, 17.7, 17.4},
  {17.7, 17.7, 16.7},
  {15.6, 16.3, 15.8},
  {15.2, 15.9, 15},
  {14.7, 15.4, 14.8},
  {14, 14.3, 14.3},
  {12.7, 13.8, 13.4},
  {13.2, 13.6, 12.5},
  {16.7, 13.8, 12.5},
  {18.4, 14.9, 15},
  {18.1, 17.8, 18.3},
  {19.2, 20.5, 21.6},
  {19.9, 21, 24},
  {21.3, 23, 25.7},
  {22.1, 24.9, 25.8},
  {20.4, 24.7, 24.6},
  {20.6, 24.5, 24.4},
  {20.4, 23.6, 24.5},
  {20.6, 22.6, 24.5},
  {20.3, 21.8, 23.2},
  {13.9, 22, 19},
  {9.6, 20.3, 17.5},
  {10.3, 17.5, 16.5},
  {11, 16.2, 15.4},
  {11.5, 16.6, 14.9},
  {11.2, 14.8, 14.7},
  {11.3, 13.5, 14.8},
  {10.6, 12.5, 13.9},
  {9.8, 11.7, 13},
  {9.6, 11.4, 12.4},
  {10.1, 11, 12.4},
  {10.3, 11.5, 12.6},
  {13.4, 11.7, 12.8},
  {15.3, 12.6, 13},
  {16.4, 14.1, 14.1},
  {17.1, 17.2, 16.7},
  {18.1, 18.8, 20.2},
  {19.2, 20.8, 22.5},
  {19.8, 22, 23.4},
  {20.2, 22.6, 23.5},
  {20, 22.4, 22.7},
  {18.4, 21, 22.7},
  {17.7, 20.4, 21.9},
  {17.5, 20.4, 21.5},
  {17.3, 19.8, 21.6},
  {16.5, 17.2, 20.4},
  {16.4, 13.9, 18.8},
  {15.8, 13.5, 17.4},
  {15.1, 13.2, 16.4},
  {13.9, 12.8, 15.5},
  {13.2, 12.3, 14.5},
  {12.4, 12.4, 13.6},
  {12.5, 12, 13},
  {12.2, 11.9, 12.9},
  {12, 11.8, 12.7},
  {13.1, 11.8, 12.8},
  {13.9, 12.7, 13.6},
  {14.2, 13.8, 14.8},
  {15.4, 15, 17},
  {16.3, 16.2, 19.2},
  {18.1, 17.7, 20.6},
  {18.5, 19.3, 21.9},
  {18.9, 21.3, 23.4},
  {18.1, 22.4, 23.7},
  {18.8, 21.6, 22.9},
  {19.2, 21.7, 22.6},
  {20, 20.9, 22.5},
  {19.3, 20.8, 22.5},
  {18.4, 21.1, 22.4},
  {18.1, 19.8, 21.3},
  {17, 18.8, 18.9},
  {16.8, 18.5, 17.9},
  {16, 18.2, 17.6},
  {15.9, 18, 17.3},
  {16.3, 18.1, 16.8},
  {16.7, 17.5, 16.1},
  {15.5, 17.7, 15.4},
  {15, 17.5, 15.1},
  {15.4, 16.9, 15},
  {15.8, 16.8, 15.5},
  {16.3, 17.4, 16.1},
  {17.1, 18.2, 17.3},
  {17.9, 18.6, 18.8},
  {19.4, 19.3, 20.4},
  {20, 20.7, 22.2},
  {20.1, 22.4, 22.9},
  {21.6, 23, 25},
  {22.1, 24.5, 26.4},
  {22.4, 24.6, 26.3},
  {21.7, 24.5, 25.7},
  {21.2, 24.4, 25.4},
  {20.8, 23.4, 25.1},
  {20.4, 22.6, 24.5},
  {19.5, 21.8, 23},
  {19.5, 21.6, 20.7},
  {19, 20.5, 19.8},
  {19.4, 20.1, 19.1},
  {18.9, 20.1, 18.4},
  {18.5, 19.7, 18.4},
  {18.3, 19.3, 18.1},
  {17.5, 19.3, 17.5},
  {17.8, 19.2, 16.9},
  {17.9, 19.6, 16.7},
  {18, 18.8, 16.7},
  {18.9, 19.4, 17.4},
  {19.3, 20, 18.6},
  {20.9, 20.6, 20.8},
  {22.1, 22.5, 23.1},
  {22.8, 23.9, 25.4},
  {23.3, 25.2, 27.2},
  {23.7, 26.2, 27.4},
  {23.9, 26.8, 26.9},
  {23.5, 26.4, 26.6},
  {22.7, 24.7, 26.9},
  {22.1, 24.6, 26.6},
  {22, 24.4, 26.7},
  {21.2, 23.8, 25.5},
  {19.9, 23.2, 24.9},
  {18.4, 21.8, 22.6},
  {18.7, 21.4, 20.8},
  {19.4, 20.8, 19.4},
  {19.1, 20.2, 18.5},
  {18, 20.5, 17.8},
  {17.2, 20.5, 17.5},
  {16.8, 20.1, 17.6},
  {16.5, 19.3, 17.3},
  {16.5, 18.7, 17},
  {17.4, 18.5, 16.5},
  {19, 19.5, 17.1},
  {20.3, 20.4, 18.5},
  {21.6, 21.8, 21.2},
  {22.2, 23, 24.1},
  {23.5, 24.2, 26.4},
  {24.5, 25.8, 28.3},
  {25.4, 27.8, 29.2},
  {25.8, 28.7, 28.9},
  {25.7, 28.9, 28.7},
  {24.9, 28.3, 29.3},
  {24.1, 27.8, 28.3},
  {23.4, 26.9, 27.8},
  {21.9, 26.1, 27.1},
  {20.2, 24.4, 25.5},
  {19.6, 23.4, 22.2},
  {19.4, 22.7, 20.4},
  {18.5, 22, 19.7},
  {18, 21.6, 18.9},
  {17.8, 20.7, 18},
  {17.6, 20.1, 17.6},
  {17.5, 19.3, 17},
  {17, 18.8, 16.5},
  {17.3, 18.5, 16.2},
  {17.1, 18.7, 16},
  {19.9, 19, 16.6},
  {22, 19.9, 19},
  {22.1, 21.5, 22.4},
  {22.8, 22.9, 24.4},
  {24.6, 24.9, 27.1},
  {25.5, 26.9, 29.3},
  {26.6, 28.9, 30.4},
  {27.1, 29.7, 30},
  {27.4, 30, 29.9},
  {26.1, 29.7, 30},
  {25.6, 29.2, 29.5},
  {25.1, 28.2, 29.4},
  {23.9, 27.2, 28.4},
  {23.3, 25.9, 26.6},
  {22.6, 24.8, 23.5},
  {20.1, 24.3, 21.4},
  {20, 23.2, 20.4},
  {19.9, 22.3, 19.4},
  {19, 21.9, 18.7},
  {18.5, 20.8, 18},
  {18.5, 20, 17.6},
  {18, 19.7, 17},
  {17.5, 19.6, 16.5},
  {17.9, 19.7, 16.2},
  {20.5, 20.2, 16.9},
  {23, 21, 19.1},
  {23.8, 23, 22.1},
  {24.8, 24.2, 25.1},
  {25.7, 26.1, 27.9},
  {26.9, 28.4, 30.2},
  {27.9, 29.9, 30.7},
  {27.6, 30.5, 30.9},
  {27.3, 30, 30.6},
  {26.6, 29.4, 30.7},
  {26.6, 29.2, 29.8},
  {26.1, 29.9, 30.2},
  {24.1, 28.7, 29.3},
  {23.3, 26.9, 27.5},
  {22, 24.9, 25.2},
  {22.3, 25.4, 22},
  {20.7, 25.2, 20.5},
  {20, 23.4, 19.4},
  {19.4, 22.4, 18.8},
  {19.6, 22.4, 18.5},
  {19.6, 21.7, 18.2},
  {19, 21.2, 17.9},
  {18.8, 20.9, 17.3},
  {18.9, 20.1, 16.8},
  {21.4, 20.6, 17.2},
  {24.3, 21.4, 19.7},
  {24.7, 24, 22.7},
  {25, 25.4, 25.4},
  {25.7, 26.9, 28.4},
  {26.9, 29, 30.6},
  {27.6, 30.2, 32.1},
  {27.2, 30.7, 31.8},
  {25.9, 30.7, 31.6},
  {25.5, 30.1, 30.5},
  {25.4, 29.3, 29.5},
  {24.5, 27.8, 28.4},
  {23.5, 27.2, 27.8},
  {22.9, 26.2, 27.1},
  {21.4, 24.8, 24.3},
  {20.2, 24.1, 21.9},
  {19.6, 23.8, 20.3},
  {19.4, 23.6, 19.2},
  {19.2, 22.8, 18.6},
  {19.1, 21.7, 17.9},
  {18.4, 20.9, 17.2},
  {17.9, 21.1, 16.7},
  {18, 20.9, 16.7},
  {18.3, 20.6, 16.9},
  {20.5, 20.9, 18.1},
  {21.4, 21.5, 20.4},
  {21.1, 22.1, 23.3},
  {22.3, 22.7, 25.3},
  {22.7, 24.2, 27.7},
  {22.9, 25.3, 28.7},
  {23.2, 25, 27.9},
  {23, 21.7, 28},
  {23.5, 21.3, 28.4},
  {24.3, 20.6, 28.4},
  {24.1, 19.8, 26.9},
  {21.8, 20, 26.3},
  {18.8, 19.2, 24.8},
  {18.4, 18, 24},
  {16.3, 17.3, 22.8},
  {15.7, 17.3, 20.2},
  {14.6, 17.2, 18},
  {14.3, 17, 16.6},
  {14.1, 16.4, 15.5},
  {13.7, 15.9, 14.8},
  {13.8, 15.6, 14},
  {13, 15.2, 13.3},
  {13, 15, 12.7},
  {12.7, 15.2, 12.3},
  {16.3, 15, 12.6},
  {17.4, 16.4, 14.5},
  {18.5, 18.7, 18.2},
  {19.8, 20.8, 21.9},
  {21.1, 23, 24.9},
  {22.7, 24.2, 27.6},
  {24, 25.9, 28.8},
  {24.6, 27.6, 29.3},
  {23.9, 28.3, 29.2},
  {23.8, 28.1, 28.4},
  {24, 27, 27.3},
  {23.3, 26.2, 26.9},
  {21.6, 25, 25.6},
  {20.3, 23.1, 24.5},
  {18.5, 21.8, 21},
  {17.2, 21.5, 18.1},
  {16.6, 21.4, 17.2},
  {17.5, 20.7, 16.4},
  {18.1, 20.2, 15.9},
  {19.3, 19.9, 16},
  {19.6, 19.7, 16},
  {18.8, 19.5, 16.2},
  {16.5, 19.3, 16.4},
  {16.7, 17.8, 15.7},
  {18.3, 18.8, 15.7},
  {19.7, 20, 17.6},
  {20.4, 21.6, 20.5},
  {20.5, 23.1, 22.3},
  {19.4, 23.5, 23.8},
  {20.4, 21.5, 24.2},
  {20.2, 22.1, 26.4},
  {20.2, 20.8, 23.6},
  {18.6, 21, 22.4},
  {18.2, 20.7, 21.8},
  {19.3, 20.1, 22.7},
  {18, 19.7, 22.1},
  {16.9, 19, 21.3},
  {16.1, 18.4, 20.7},
  {16.5, 18, 20.1},
  {16, 17.5, 19.4},
  {14.8, 16.6, 17.8},
  {14.4, 16.3, 16.9},
  {13.5, 16.1, 16.4},
  {13.3, 15.4, 16},
  {12.8, 14.8, 14.8},
  {11.6, 15, 14.5},
  {11.2, 15.2, 14.1},
  {11.4, 15, 13.7},
  {13.2, 14.8, 13.9},
  {15.2, 15, 14.6},
  {15.4, 15.9, 15.5},
  {16.7, 17.1, 17.9},
  {17.3, 18.9, 20.2},
  {17.7, 19.7, 22.3},
  {18.3, 20.3, 23.6},
  {19.3, 22.3, 24.5},
  {20.6, 23.4, 25.7},
  {20.7, 23.1, 24.9},
  {19.9, 21.9, 21.7},
  {18.4, 22, 21.9},
  {17.7, 22, 22.9},
  {16.6, 20.4, 20.1},
  {16.9, 19.2, 18.3},
  {16.9, 18.6, 16.7},
  {16, 18.5, 15.2},
  {16, 18.3, 14.3},
  {16.4, 18.1, 13.6},
  {16.7, 17.1, 13},
  {15.8, 17, 11.9},
  {15.6, 17, 11.2},
  {14.8, 16.3, 10.7},
  {13.3, 16, 10.2},
  {16, 16.2, 10.3},
  {18, 16.7, 13.2},
  {18.6, 18.4, 17},
  {19.7, 20.4, 20.6},
  {20.6, 21.8, 24.2},
  {21.3, 22.7, 25.5},
  {20.7, 23.2, 25.7},
  {19, 23.3, 24.8},
  {19.4, 23.4, 25.3},
  {20, 23.3, 25},
  {19.9, 22.8, 24.6},
  {19.2, 22, 24.7},
  {17, 20.9, 24.4},
  {16.5, 18.9, 22.8},
  {16, 17.6, 21},
  {15, 16.9, 17.6},
  {14.1, 16.4, 15.6},
  {14.1, 15.8, 13.1},
  {13.7, 15.2, 11.3},
  {13.2, 14.8, 9.7},
  {11.9, 13.8, 8.8},
  {11.1, 13, 8.2},
  {9.3, 12.6, 7.4},
  {9.4, 12.3, 6.9},
  {13, 12.5, 6.9},
  {15.2, 13.1, 9.6},
  {15.8, 15.5, 14},
  {16.8, 18.1, 18.1},
  {18.1, 20.1, 21.2},
  {19.3, 22.1, 23.3},
  {20.4, 23.1, 24.5},
  {21.8, 24.3, 25.5},
  {21.9, 25.2, 26.5},
  {20.5, 25.6, 26.1},
  {20, 25.5, 24.3},
  {18.6, 23.7, 24},
  {17.4, 22.2, 22.5},
  {15.8, 19.9, 19.1},
  {15.9, 18.9, 15.7},
  {15.6, 18.1, 13.8},
  {14.8, 16.9, 13},
  {13.6, 15.8, 12.1},
  {12.6, 15.1, 11.4},
  {12.6, 15, 10.7},
  {11.7, 13.8, 10.3},
  {11.4, 13.6, 10},
  {11.1, 13.3, 9.8},
  {11.7, 13.5, 9.8},
  {14.9, 14.1, 10.8},
  {17.4, 15.3, 13.3},
  {17.5, 16.6, 16.1},
  {18.9, 18.6, 19.4},
  {19.1, 19.9, 21.8},
  {20.1, 21.4, 23.8},
  {21, 23.1, 25.3},
  {20.9, 24.2, 24.9},
  {20.1, 23.9, 24},
  {19.1, 22.4, 22.6},
  {18, 21.3, 22.5},
  {17.4, 20.3, 21.9},
  {16.6, 19.7, 21.2},
  {15.9, 18.8, 20.5},
  {14.4, 18, 18.4},
  {14.5, 17.7, 17.4},
  {14.4, 17.3, 16.8},
  {14.3, 16.7, 16.3},
  {13.6, 16.5, 15.7},
  {13.8, 16.2, 15.2},
  {13.7, 14.2, 14.9},
  {13.2, 13.5, 14.8},
  {13.1, 13.2, 14.7},
  {14, 13, 14.6},
  {14.3, 13.6, 14.7},
  {14.3, 15.4, 15.3},
  {14.2, 17.2, 16.1},
  {14.9, 17.3, 17.3},
  {16.2, 18.1, 20.4},
  {16.2, 18.8, 20.2},
  {16.5, 16.6, 18.8},
  {14.6, 18.3, 17.5},
  {14.4, 18.8, 17.8},
  {12.6, 18, 16.8},
  {12.2, 17.5, 16.4},
  {12.2, 17.1, 16.6},
  {11.7, 16.2, 16.4},
  {10.8, 14.4, 14.2},
  {11.6, 12.7, 12.7},
  {10.7, 12.7, 12.2},
  {9.2, 12.8, 12.1},
  {7.9, 12.7, 11.5},
  {7.3, 11.8, 10.4},
  {6.8, 11.8, 9.2},
  {6.8, 10.8, 8.6},
  {6.4, 9.7, 7.6},
  {5.9, 9.4, 6.9},
  {5.9, 9.2, 6.3},
  {8.9, 9.6, 6.2},
  {12, 10.6, 8},
  {12.9, 13.3, 11.4},
  {14, 15.8, 15.1},
  {15.1, 17.2, 18.3},
  {16.6, 18.8, 20.9},
  {17.2, 20, 21.9},
  {17.8, 21.2, 22.8},
  {17.5, 21.5, 23.3},
  {17.3, 21.7, 22.8},
  {17.2, 21.2, 21.4},
  {16.3, 19.6, 19.6},
  {15, 17.8, 18.2},
  {13.2, 16.3, 16.3},
  {11.8, 15.7, 12.7},
  {10.7, 15.3, 11.7},
  {10.2, 14.7, 10.5},
  {10.2, 13.6, 9.7},
  {11.6, 13, 9.1},
  {11.9, 12.9, 8.5},
  {11.2, 13.3, 8.7},
  {9.1, 12.5, 8.9},
  {9, 11.4, 8.1},
  {9.2, 11.9, 7.9},
  {10.9, 12.3, 8.4},
  {13.2, 12.8, 9.8},
  {14.6, 14.1, 12.5},
  {16.2, 15.7, 15.4},
  {16.9, 17.9, 19.2},
  {17.8, 19.4, 21.2},
  {17.7, 20.7, 22.2},
  {17.9, 21.5, 22.7},
  {18.4, 21.8, 23},
  {18.6, 22, 23},
  {19.1, 21.9, 22.8},
  {18.6, 21.4, 22.4},
  {17.4, 20.3, 21.5},
  {14, 18.2, 19.1},
  {12.6, 16.8, 16.1},
  {13.7, 16.8, 13},
  {14.6, 16.2, 12},
  {13.7, 15.7, 11.1},
  {14.1, 15.3, 10.1},
  {13.6, 14.9, 9.7},
  {11.5, 13.6, 9.2},
  {10.7, 12.6, 8.6},
  {10.3, 11.6, 8.2},
  {10.6, 11.4, 8.2},
  {12.6, 11.8, 8.4},
  {15.4, 13.2, 10.4},
  {17, 15.7, 14.3},
  {18.1, 17.5, 17.9},
  {19, 19.8, 20.9},
  {20, 21.5, 23.1},
  {21, 22.8, 24.1},
  {19.5, 23.7, 24.1},
  {19.6, 23, 23},
  {19.3, 22.3, 22.9},
  {19.5, 21.5, 22.5},
  {18.4, 21, 22.7},
  {17.1, 20, 21.9},
  {16.1, 18.4, 20.2},
  {14.1, 17.4, 17.5},
  {13.6, 16.8, 15.6},
  {13.8, 16.4, 14.5},
  {14.1, 16.1, 13.3},
  {13.6, 16.5, 12.8},
  {13.3, 16.3, 12.4},
  {13.2, 16.1, 12.2},
  {14.3, 14.9, 12},
  {13.8, 15, 12},
  {13.6, 14.6, 11.9},
  {15.1, 15.8, 12.7},
  {16.6, 16.3, 14.8},
  {17.5, 17.3, 18},
  {17.4, 18.4, 20.8},
  {17.9, 20.1, 21.6},
  {18.5, 21.2, 23.2},
  {18.1, 21.8, 22.7},
  {18, 21.5, 22.1},
  {19.8, 22.1, 23.5},
  {19.1, 22.1, 23.5},
  {18.7, 21.6, 22.5},
  {18.3, 19.4, 20.8},
  {17.5, 17.7, 21.2},
  {15.8, 17, 20.4},
  {15.7, 16.7, 19.1},
  {15.9, 16.2, 18.3},
  {15.8, 15.9, 17.5},
  {15.3, 15.2, 17.2},
  {15.1, 15, 16.8},
  {14.6, 15.1, 16.4},
  {12.8, 15.3, 16.3},
  {12.2, 15.1, 16},
  {12, 14.5, 15.7},
  {12, 14.2, 15.5},
  {13, 14.2, 15.6},
  {13.9, 14.8, 16},
  {15.7, 15.5, 16.8},
  {17.4, 16.6, 18.6},
  {18.4, 18.4, 21.5},
  {19.3, 21.7, 23.6},
  {20.1, 22.6, 24.6},
  {20.1, 23.4, 23.3},
  {20.1, 23.7, 23.5},
  {20, 23.1, 23.3},
  {19.5, 22.6, 23.5},
  {18.2, 21.6, 22.6},
  {17.9, 20.4, 22.2},
  {17.3, 18.8, 21.2},
  {16.9, 18.1, 19.4},
  {16.6, 17.6, 18},
  {16.1, 17.8, 16.9},
  {16, 16.3, 15.9},
  {14.9, 16.1, 15.6},
  {15.1, 15.8, 15.1},
  {14.4, 15.3, 14.9},
  {13.4, 15.2, 14.3},
  {12.9, 15.1, 13.6},
  {12.8, 14.9, 12.8},
  {13.7, 14.7, 12.8},
  {16.3, 15.6, 14.3},
  {17.2, 17.9, 16.9},
  {17.7, 18.5, 20.4},
  {19.9, 19.9, 23},
  {21.3, 20.7, 24.6},
  {21.1, 23.1, 25},
  {19.9, 22.2, 23.7},
  {18, 21.5, 21},
  {17.5, 21, 21.6},
  {16.7, 20.7, 20.7},
  {15.9, 20, 20.9},
  {15.7, 18.9, 19.7},
  {15.6, 16.5, 18.7},
  {16.1, 15.6, 17.5},
  {15.7, 14.2, 16.9},
  {14.7, 13.6, 16.6},
  {13.4, 13, 15.7},
  {12.8, 12.5, 15.2},
  {12.5, 12.4, 14.3},
  {12.9, 12.2, 13.8},
  {12.9, 11.9, 13.1},
  {12.7, 11.7, 12.4},
  {13.5, 11.4, 12.1},
  {13.7, 11.9, 12.8},
  {13.9, 12.5, 13.9},
  {14.5, 13.9, 15},
  {15.4, 15.2, 17.4},
  {16.8, 16.7, 19.7},
  {17.3, 18, 20.7},
  {17.7, 19.4, 21.4},
  {16.3, 19.2, 20.3},
  {15.1, 17.9, 19.3},
  {15, 17, 18.9},
  {15, 16.6, 18.7},
  {14.7, 15.8, 17.6},
  {14.1, 15.5, 17.3},
  {13.1, 15, 17},
  {12.3, 14.3, 16.5},
  {11.6, 14.1, 15.3},
  {11.3, 13.6, 14.9},
  {11.1, 13.1, _},
  {11, 12.9, _},
  {10.7, 12.7, _},
  {10.1, 11.9, _},
  {9.8, 11.9, _},
  {9.9, 11.5, _},
  {10, 11.7, _},
  {10.1, 11, _},
  {12.9, 12, _},
  {14.1, 14.1, _},
  {14.8, 16.5, _},
  {16.9, 18.3, _},
  {18.5, 19.7, _},
  {17.9, 20.5, _},
  {18.8, 20, _},
  {18.5, 20, _},
  {19, 20.5, _},
  {18.9, 20.7, _},
  {17.8, 19.9, _},
  {15.1, 19, _},
  {13.2, 16.6, _},
  {11.3, 15.3, _},
  {10.6, 14.7, _},
  {10.2, 14.8, _},
  {10.2, 14.1, _},
  {9.5, 13.2, _},
  {9.8, 13, _},
  {9.1, 12.4, _},
  {9.6, 12.4, _},
  {10.4, 11.8, _},
  {10.3, 11.4, _},
  {11.3, 11.5, _},
  {13.2, 13.3, _},
  {14.6, 15.4, _},
  {15.9, 17.1, _},
  {16.8, 19.4, 16.9},
  {18.9, 20.4, 20.8},
  {20.5, 21.7, 24},
  {20.8, 22.5, 25.4},
  {21.8, 22.1, 25.8},
  {22, 22.4, 25.3},
  {20.9, 21.9, 25.5},
  {19, 21.4, 24.4},
  {17.1, 19.8, 23.3},
  {15.1, 18.5, 19.7},
  {12.8, 17.8, 15.7},
  {12.4, 17.1, 14.2},
  {12.4, 15.6, 12.8},
  {12.4, 14.8, 11.5},
  {11.8, 14.3, 10.8},
  {11.1, 14.2, 9.8},
  {10.1, 13.6, 9.1},
  {10.4, 13.3, 8.7},
  {10.7, 13.1, 8.2},
  {10.5, 12.7, 7.8},
  {12, 12.7, 7.9},
  {15.4, 13.6, 11.2},
  {17.3, 16, 15},
  {18.3, 18.4, 19.2},
  {19.5, 20.5, 22},
  {20.7, 23.3, 24.3},
  {22.3, 24.9, 26.5},
  {23.6, 25.6, 27.8},
  {23.7, 26.9, 27.2},
  {23.9, 26.5, 26.1},
  {23.5, 26.2, 26},
  {21, 25.1, 24.8},
  {19.2, 23.3, 22.9},
  {16.3, 21.4, 18.8},
  {16.2, 20.4, 16.2},
  {15, 20.2, 14.8},
  {15, 19.7, 14.2},
  {14.2, 18.6, 13.4},
  {14.5, 18.3, 12.9},
  {13.6, 17.8, 12.3},
  {13.1, 16, 11.8},
  {12.7, 15.2, 11.3},
  {12.7, 14.3, 10.6},
  {12.5, 13.9, 10.6},
  {13.7, 14.3, 11.4},
  {17.4, 15.3, 13.3},
  {19.2, 17, 17.8},
  {19.8, 20.1, 20.9},
  {20.3, 21.7, 23.6},
  {21.4, 23.1, 25.2},
  {21.7, 24.2, 25.3},
  {21.5, 24.9, 25.1},
  {21.4, 25, 25},
  {21, 24.7, 25},
  {20.5, 23.4, 24.1},
  {19.3, 21.8, 23.2},
  {18.8, 21, 22.7},
  {18.1, 19.8, 21.5},
  {17.8, 19.9, 19.8},
  {16.6, 19.6, 18.3},
  {16.6, 18.5, 17.1},
  {15.9, 16.3, 16.8},
  {15.9, 15.2, 16.8},
  {15.9, 15.5, 17.1},
  {14.6, 14.4, 16.6},
  {13.4, 14.1, 15.3},
  {13.3, 13.9, 14.6},
  {13.8, 13.8, 14.3},
  {14.5, 14.4, 14.3},
  {16.1, 14.8, 16.9},
  {17.1, 17.3, 19.9},
  {18.2, 19.3, 22},
  {20.1, 20.9, 24.2},
  {21.5, 22, 25.9},
  {22.4, 24, 25.9},
  {22.6, 24.5, 24.5},
  {20.4, 23.2, 24},
  {19.2, 22.6, 24.2},
  {18.8, 22.3, 23.5},
  {18.8, 21.8, 22.6},
  {17.4, 20.8, 21.5},
  {15.5, 19.2, 19.8},
  {15.1, 18.1, 17.2},
  {15.1, 17.8, 15.9},
  {14.8, 17.2, 15.1},
  {15.4, 16.7, 14.4},
  {15.2, 16.5, 13.8},
  {14.5, 16.4, 13.5},
  {14.8, 16.1, 13.3},
  {15.4, 16, 13.3},
  {15.3, 16.1, 13.1},
  {14.8, 16.1, 12.9},
  {15.6, 16.8, 13.7},
  {15.3, 16.8, 14.7},
  {15, 16.6, 14.8},
  {15.1, 15.6, 15.3},
  {15.6, 14.8, 15.6},
  {14.7, 13.3, 15.8},
  {14.4, 12.7, 16},
  {13.7, 12.4, 15.9},
  {13.7, 12.4, 16},
  {13.8, 14.2, 18.2},
  {13.8, 15, 18.8},
  {13.7, 15.3, 18.6},
  {12.9, 14, 17.4},
  {11.8, 12.9, 15.4},
  {12, 12.9, 14.1},
  {12.1, 12.7, 13.5},
  {11.6, 12.9, 13},
  {11.3, 13, 12.6},
  {11.3, 13, 12.5},
  {11.8, 12.9, 12.7},
  {11.9, 12.8, 12.8},
  {11.8, 12.5, 12.9},
  {11.7, 12.2, 12.9},
  {11.5, 11.9, 12.9},
  {11.4, 11.7, 13},
  {11.2, 11.8, 13.2},
  {11.5, 11.9, 13.4},
  {11.4, 12, 13.7},
  {11.3, 12.3, 13.8},
  {11.4, 12.8, 14.2},
  {11.6, 13, 14.5},
  {11.8, 13.4, 14.9},
  {12.3, 13.4, 15.2},
  {12.5, 13.4, 15.3},
  {12.8, 13.3, 15.7},
  {12.9, 13.3, 15.8},
  {12.3, 12.9, 15.7},
  {11.9, 12.2, 14.6},
  {12.3, 12.5, 14},
  {12.2, 12.1, 13.7},
  {11.9, 12.3, 13.1},
  {11.3, 12.5, 13.4},
  {10, 12, 13.2},
  {9.4, 11.7, 12.5},
  {9.5, 12.2, 12.2},
  {9.3, 12.4, 12.2},
  {9, 12.4, 12},
  {9.9, 12.5, 12},
  {10.6, 12.5, 12.4},
  {11.5, 12.5, 12.8},
  {12.4, 12.5, 13.2},
  {12.5, 12.6, 13.7},
  {12.3, 13.2, 14.2},
  {12.5, 13.1, 14.8},
  {12.3, 13.8, 15.7},
  {12.6, 13.3, 16},
  {12.7, 13.6, 15.3},
  {12.7, 13.8, 15},
  {13, 13.8, 15.2},
  {12.8, 13.7, 15.4},
  {12.3, 13.4, 15.2},
  {11.8, 13.1, 14.8},
  {11.6, 12.7, 14.6},
  {11.4, 12.5, 14.4},
  {11.2, 12.6, 14.2},
  {11.1, 12.7, 14},
  {11.1, 12.6, 13.7},
  {11.2, 12.5, 13.6},
  {11.1, 12.5, 13.6},
  {11, 12.3, 13.4},
  {10.8, 12.1, 13.2},
  {10.7, 11.7, 13.2},
  {11.2, 12.1, 13.3},
  {11.4, 12.7, 13.4},
  {11.7, 13, 13.5},
  {12.6, 14.1, 14},
  {14.2, 15.2, 15.2},
  {15.8, 17, 17.5},
  {16.6, 18.9, 19.2},
  {16.5, 19.5, 19.8},
  {17, 19.5, 20.2},
  {17.6, 18.9, 21.3},
  {17.2, 18.9, 21},
  {17.2, 19.1, 20.3},
  {14.8, 18.4, 18.5},
  {13.7, 15.9, 16.5},
  {13.9, 15.1, 15.3},
  {13.7, 15, 14.6},
  {13.1, 14.8, 14.2},
  {12.6, 14.9, 13.9},
  {12.3, 14.7, 13.6},
  {12.6, 14.1, 13.6},
  {11.7, 13.7, 12.8},
  {11.7, 13.4, 12.2},
  {11.8, 13.3, 12.2},
  {11.1, 12.5, 12.5},
  {11.8, 12.2, 12.8},
  {14.2, 13.2, 13},
  {15.5, 14.8, 15.1},
  {17.2, 17.3, 18.3},
  {18.3, 19.6, 21.3},
  {19.5, 21.1, 23.7},
  {20.1, 21.1, 25},
  {20.7, 22.6, 24.6},
  {20.9, 23.5, 23.7},
  {21, 23.2, 23.7},
  {20.8, 22.7, 23.4},
  {18.2, 21.7, 21.8},
  {16.9, 19.6, 19.5},
  {15.9, 18.1, 17.2},
  {15.2, 17.7, 15.6},
  {15.9, 17, 15.1},
  {15.3, 17.2, 15.1},
  {15.5, 17.4, 15.3},
  {13.8, 16.2, 14.6},
  {13.4, 15.8, 14},
  {13.4, 15.7, 13.4},
  {12.8, 15.3, 13.2},
  {13.2, 15, 13.2},
  {14, 15.2, 13.6},
  {14.4, 15.1, 14.1},
  {15.1, 15.8, 15.3},
  {16, 16.2, 16.9},
  {17, 17.3, 19.1},
  {17.9, 19, 20.8},
  {18.8, 20.1, 22.2},
  {19.2, 21.1, 21.9},
  {17.2, 20.2, 20.9},
  {17.4, 19.5, 21.5},
  {17.6, 19.3, 22},
  {16.9, 19.3, 21.7},
  {17.4, 19.2, 21.5},
  {17.1, 18.8, 20.7},
  {16.6, 18.1, 19.4},
  {16.7, 18, 18.3},
  {16.7, 17.7, 17.4},
  {16.5, 17.8, 16.7},
  {15, 18.1, 16.5},
  {14.3, 17.5, 16.5},
  {13.9, 17.3, 16.3},
  {13.7, 16.6, 15.8},
  {14, 15.8, 14.9},
  {13.4, 16.2, 14.1},
  {13.2, 16.3, 14.2},
  {14.2, 16.2, 14.5},
  {16.4, 16.9, 15.9},
  {17.2, 17.8, 17.6},
  {17.4, 18.7, 19.6},
  {18.2, 19.5, 22.1},
  {19.3, 21, 23},
  {20.2, 22.1, 23.4},
  {19.6, 22.7, 23.6},
  {20, 22.4, 23.5},
  {19.2, 22.2, 22.8},
  {18.5, 21.9, 22.6},
  {18.5, 21, 22.1},
  {18, 19.9, 21.2},
  {17.5, 19.5, 20.3},
  {16.8, 18.6, 18.9},
  {16.2, 18.2, 18.4},
  {15.5, 18, 18.1},
  {15.1, 18, 17.2},
  {16.1, 17.4, 16.9},
  {15.6, 17.5, 16.6},
  {15.3, 17.4, 16.7},
  {15.2, 16.9, 16.8},
  {15.4, 16.6, 16.6},
  {15, 16.3, 16.5},
  {15.3, 16.5, 16.5},
  {16.1, 16.8, 17.1},
  {16.3, 17.8, 19.2},
  {17.2, 18.4, 21.8},
  {18.7, 19.5, 22.6},
  {19.1, 20.6, 22.2},
  {19.5, 21.5, 23.2},
  {19.1, 22.2, 22.7},
  {18.3, 21.3, 22.5},
  {17.7, 20.7, 22.8},
  {17.4, 19.9, 21.8},
  {17.4, 19.4, 21},
  {16.4, 18.8, 20.3},
  {15.6, 17.5, 18.9},
  {15.1, 15.4, 17.6},
  {14.8, 14.5, 16.7},
  {14.5, 13.9, 16.3},
  {14.1, 13.8, 16.2},
  {14.1, 13.8, 16.1},
  {13.8, 13.9, 15.9},
  {13.6, 13.9, 15.7},
  {13.1, 13.9, 15.5},
  {12.9, 14, 15.3},
  {12.8, 13.9, 15.1},
  {12.7, 13.9, 15.2},
  {12.8, 14.2, 15.4},
  {13.3, 15.1, 15.8},
  {13.9, 16, 16.6},
  {14.6, 16.5, 18.5},
  {15.2, 18.1, 20.8},
  {16.5, 19.5, 22.1},
  {17.6, 20.2, 23.1},
  {17.4, 20.4, 23},
  {16.8, 19.6, 22.1},
  {16.9, 18.9, 20.3},
  {16, 18, 19.7},
  {15.5, 17.2, 19.1},
  {15.1, 16.6, 18.1},
  {14.8, 16.3, 17.5},
  {14.7, 15.9, 17.3},
  {14.7, 15.9, 16.3},
  {14.8, 15.9, 16},
  {15, 15.8, 16.1},
  {13.9, 15.2, 15.9},
  {13.7, 14.8, 15.2},
  {14, 14.7, 14.5},
  {14, 14.2, 13.7},
  {14.1, 14.3, 13.2},
  {14.3, 14.3, 13.6},
  {15.8, 14.6, 14.6},
  {17.9, 16.3, 17.4},
  {18.8, 18.4, 20.6},
  {20.1, 20, 23.2},
  {20.8, 21.5, 25.3},
  {21.5, 22.8, 26.2},
  {22.1, 24, 25.2},
  {22.6, 24.7, 24.8},
  {22.2, 24.6, 24.1},
  {21.9, 23.9, 24.1},
  {19.8, 23, 23.8},
  {17.8, 21.1, 21.2},
  {16.8, 19.8, 18.8},
  {16.3, 19.2, 17.4},
  {15.8, 17.7, 16.5},
  {14.9, 17.4, 15.7},
  {14.6, 16.9, 15.1},
  {14.5, 16.2, 14.6},
  {14.3, 16.1, 14.2},
  {14.6, 15.8, 13.8},
  {14.3, 15.4, 13.4},
  {14.4, 15.5, 13.1},
  {13.8, 14.8, 13.6},
  {14.1, 15.1, 14.3},
  {16.5, 16, 15},
  {18.9, 17.5, 16.4},
  {19.9, 20.4, 20.3},
  {21.2, 21.2, 23.4},
  {22.3, 22.2, 25.6},
  {23.1, 23.9, 27.6},
  {23.8, 25.4, 27.8},
  {24, 26.4, 26.8},
  {23.6, 26.2, 26.4},
  {22.6, 25.5, 25.9},
  {21.5, 24.3, 24.4},
  {19.8, 22.3, 22.5},
  {18.5, 21.1, 20.2},
  {18.4, 20.8, 19},
  {18.7, 20.3, 18.4},
  {18.5, 19.4, 18.1},
  {17.7, 19, 17.9},
  {16.6, 18.4, 17.6},
  {16.3, 18.7, 17.6},
  {16.7, 18.5, 17.8},
  {16.7, 18.3, 17.9},
  {17.2, 17.7, 18},
  {17.2, 17.4, 18.1},
  {17.3, 18, 18.3},
  {18, 18.8, 19},
  {18.5, 19.6, 20.6},
  {19.3, 20.3, 22.8},
  {19.5, 21.2, 23.6},
  {20.9, 22.9, 25.2},
  {22, 24, 25.7},
  {22.6, 24.5, 25.5},
  {22.1, 24.4, 25.3},
  {20.7, 24.2, 25.1},
  {20.2, 23.5, 24.4},
  {19.6, 22.4, 23.8},
  {18.7, 20.9, 22.6},
  {17.3, 19.8, 21.3},
  {16.3, 19.5, 20.7},
  {16.2, 19.5, 20},
  {16.3, 19.4, 19.4},
  {16.9, 19.2, 19.2},
  {16.3, 19.5, 19.1},
  {16.1, 18.9, 18.8},
  {16.6, 18.5, 18.5},
  {16.8, 17.7, 18.1},
  {16, 16.7, 17.8},
  {15.9, 16.5, 17.5},
  {16.5, 17, 17.2},
  {17.6, 18.1, 18},
  {18.5, 19.5, 19},
  {19.7, 20.1, 20.7},
  {20.4, 21, 22.8},
  {21.7, 22.6, 24.7},
  {23.1, 24.2, 26},
  {23.4, 25.6, 26.7},
  {24.1, 25.5, 27.6},
  {23.4, 25.5, 26.2},
  {22, 24.2, 24.5},
  {20.8, 23.6, 24.3},
  {19.4, 21.9, 22.8},
  {17.3, 20.6, 20.4},
  {17.4, 20.2, 19.2},
  {17.2, 19.5, 18.9},
  {17.4, 19, 18.6},
  {16.9, 18.4, 17.9},
  {17, 18.2, 17.6},
  {17, 18.6, 17.5},
  {16.5, 18.4, 17.4},
  {16.5, 17.8, 16.7},
  {15.5, 17.5, 15.9},
  {15.5, 17.3, 15.4},
  {15.8, 17.3, 15.5},
  {18, 18, 16.7},
  {20.5, 19.5, 18.8},
  {21.1, 21.6, 22.6},
  {22.7, 23.1, 25.6},
  {23.6, 25.6, 27.4},
  {24.7, 25.8, 29.3},
  {25.7, 27, 29.4},
  {23, 27.4, 28.2},
  {21.8, 24.5, 25.5},
  {21, 24.3, 22},
  {20.2, 23.8, 19.9},
  {18.6, 21.9, 19},
  {19.1, 17, 18.5},
  {18.8, 16.1, 18.4},
  {18, 15.6, 18},
  {16.9, 15.7, 17.6},
  {17.3, 15.7, 17.4},
  {16, 16, 17},
  {15.1, 15.6, 16.3},
  {14.9, 15.1, 15.7},
  {15, 15.3, 15.3},
  {14.2, 15.1, 14.8},
  {13.2, 15.1, 14.1},
  {14.6, 15.3, 13.9},
  {16.6, 16, 14.7},
  {18.8, 16.5, 16.5},
  {19.2, 18.3, 19.5},
  {20.6, 20, 22.6},
  {22.1, 22.1, 25.4},
  {22.9, 23.7, 26.7},
  {23.5, 25.4, 27.4},
  {22.9, 25.5, 25.2},
  {21.1, 23.8, 23.7},
  {19.4, 22.4, 21.9},
  {18.3, 22.4, 20.8},
  {16.7, 20.8, 19.7},
  {16.2, 19.7, 18.5},
  {15.9, 19, 17.3},
  {15.7, 16.8, 16.7},
  {16, 14.2, 16.7},
  {15.4, 13.3, 16.3},
  {13.8, 12.7, 15},
  {13, 12.5, 14.1},
  {12.6, 12.6, 13.1},
  {12.5, 12.4, 12.8},
  {12.4, 12.4, 12.5},
  {12.2, 12, 13},
  {12.2, 12, 13.5},
  {13.8, 12.7, 13.9},
  {16.2, 14.3, 14.2},
  {16.5, 16.4, 16.5},
  {18.8, 17.2, 20.4},
  {19.8, 19, 22.9},
  {20.6, 21.4, 24.4},
  {21.2, 22.6, 24.3},
  {20.8, 23.1, 24.3},
  {19.8, 23, 24.3},
  {19, 21.8, 23.4},
  {17.3, 19.9, 21.4},
  {17, 19.3, 19.5},
  {16, 18.1, 18.2},
  {14.8, 16.2, 17.2},
  {13.7, 14.1, 16},
  {13, 13.6, 15.4},
  {13, 13, 14.9},
  {12.7, 12.6, 14.5},
  {12.1, 12.3, 14.1},
  {11.6, 11.8, 13.8},
  {11.5, 11.3, 13.7},
  {11.3, 11.1, 13.6},
  {12, 10.9, 13.7},
  {12.5, 11.3, 13.9},
  {13, 12.8, 14.2},
  {14, 13.6, 14.5},
  {14.9, 14.7, 15.5},
  {16, 16.4, 18.3},
  {16.3, 18.2, 19.9},
  {16.8, 19.7, 21.2},
  {17.7, 20.5, 21.1},
  {18.2, 20.8, 21.7},
  {18.1, 20.9, 21.6},
  {18.3, 20.7, 21.3},
  {15.8, 19.5, 19.7},
  {13.4, 17.3, 17.3},
  {12.4, 16.1, 15.2},
  {12.1, 15.5, 13.9},
  {11.6, 14.7, 13},
  {12.1, 14.2, 12.4},
  {11.5, 14.6, 11.7},
  {11.3, 14.5, 11.1},
  {11.4, 13.4, 10.6},
  {10.8, 12.9, 10.1},
  {10.3, 12.1, 9.7},
  {10.2, 11.7, 9.3},
  {10.6, 11.3, 9},
  {10.2, 11.5, 9.8},
  {12.2, 12.4, 10.7},
  {15.9, 13.9, 12.2},
  {17, 16.6, 15.7},
  {18.2, 18.3, 19.3},
  {18.6, 19.7, 21.7},
  {19.2, 21, 23.6},
  {19.7, 21.9, 24.2},
  {19.9, 22.3, 24.1},
  {19.6, 22.4, 23.1},
  {18.6, 21.7, 21.9},
  {16.8, 20.2, 20.4},
  {15.2, 18, 18.5},
  {13.4, 16.7, 15.6},
  {13.1, 16.1, 14.1},
  {12, 15.6, 13.1},
  {11.6, 14.9, 12.1},
  {11.9, 14.2, 11.8},
  {12.1, 13.7, 11.2},
  {11.9, 13.5, 10.6},
  {11.7, 12.6, 10.3},
  {12.1, 11.9, 10},
  {11.6, 11.5, 9.5},
  {11.4, 11.5, 9.2},
  {12, 11.6, 9.3},
  {13.8, 12.3, 10.4},
  {16.3, 13.7, 13.7},
  {17.8, 16.4, 17},
  {17.9, 18.1, 19.9},
  {18.8, 19.2, 22.2},
  {19.6, 20.8, 23.2},
  {20.1, 22, 24.8},
  {19.9, 22.5, 24.2},
  {19.1, 22.4, 22.6},
  {18.3, 20.8, 22.2},
  {17.8, 19.8, 21.4},
  {16.4, 18.6, 20},
  {15.5, 18.2, 19.1},
  {15.3, 17.7, 17.8},
  {14.9, 16.5, 17.1},
  {14.6, 15.9, 16.6},
  {14.7, 15.4, 16.2},
  {14.8, 15.8, 16},
  {14.6, 15.9, 15.7},
  {14.2, 15.1, 14.9},
  {13.4, 14.8, 14.4},
  {13.4, 14.8, 13.8},
  {12.8, 14.5, 13},
  {13, 14.3, 12.8},
  {14.6, 14.6, 13.6},
  {16.1, 16.2, 15.4},
  {17, 18.2, 19.1},
  {17.8, 19.4, 22.2},
  {19.1, 20.9, 23.4},
  {20.5, 22.3, 24.9},
  {20.5, 23.5, 24.1},
  {20.1, 23.4, 22.8},
  {19.9, 22.9, 23.7},
  {18.3, 22.2, 22.1},
  {18.5, 19.9, 21.5},
  {17.4, 18.9, 20.3},
  {15.6, 18.6, 18.3},
  {16.8, 18.5, 17.5},
  {16.8, 18.4, 17.3},
  {16.3, 16.8, 17.4},
  {15.4, 15.8, 17.1},
  {15, 15.5, 16.9},
  {14.9, 15.3, 16.6},
  {14.6, 15, 16.5},
  {15, 14.9, 16.3},
  {15, 14.9, 16.2},
  {14.3, 14.8, 15.9},
  {14.5, 14.9, 15.9},
  {15, 15.6, 16},
  {16, 16.1, 16.4},
  {17, 16.9, 16.9},
  {16.5, 17.5, 17.6},
  {15.9, 17.1, 18.3},
  {15.3, 16.2, 17.9},
  {14.6, 16.1, 17.3},
  {15, 16, 17.1},
  {14.9, 15.7, 17.2},
  {15.3, 15.9, 16.6},
  {15.1, 15.5, 16.4},
  {14.6, 15.5, 16.3},
  {14.1, 15.1, 16.2},
  {14, 14.9, 15.8},
  {14, 14.6, 15.6},
  {13.8, 14.6, 15.4},
  {13.3, 14.5, 15.3},
  {11.9, 14.1, 15.1},
  {11.4, 13.3, 15},
  {11.5, 13.3, 14.8},
  {11.1, 13.4, 14.6},
  {10.8, 13.5, 14.5},
  {10.8, 13.7, 14.2},
  {11.2, 14, 14.5},
  {11.9, 14.5, 14.7},
  {13.9, 14.6, 15},
  {16.2, 15, 16.5},
  {17.3, 16.2, 17.9},
  {18.4, 18, 21},
  {18.8, 18.9, 23},
  {19.2, 19.5, 23.2},
  {19.4, 19.9, 22.5},
  {17.4, 19.8, 21.5},
  {16.6, 19.9, 21.1},
  {16.1, 18.6, 19.9},
  {15, 16.1, 18.6},
  {14.8, 15.8, 17.5},
  {15, 15.9, 16.8},
  {15.1, 15.8, 16.7},
  {14.7, 15.6, 16.7},
  {14, 15.5, 16.7},
  {14.3, 15.4, 16.2},
  {13.6, 15.5, 15.9},
  {13.3, 15.5, 15.8},
  {13.7, 15.2, 15.9},
  {13.4, 15.1, 16},
  {13.9, 14.9, 15.9},
  {14.4, 15.4, 16.1},
  {14.9, 16.5, 16.4},
  {15.9, 16.5, 17.5},
  {16.5, 17.8, 18.9},
  {16.5, 18.4, 18.6},
  {16.4, 16.7, 17.9},
  {16.4, 16.7, 19.6},
  {17.6, 18.7, 21},
  {17.6, 19, 20.9},
  {18.2, 19.7, 20.8},
  {18.8, 18.8, 21.8},
  {16.9, 19.1, 19.3},
  {15, 16.1, 17.9},
  {13.7, 17, 16.5},
  {13.8, 15, 15.8},
  {13.2, 14.2, 15.4},
  {12.1, 14.4, 14.3},
  {11.2, 13, 12.7},
  {10.6, 12.3, 11.8},
  {10.1, 12, 11.6},
  {10, 11.8, 11.8},
  {10.4, 11.9, 12},
  {11, 12.1, 12.1},
  {11.3, 11.9, 12.2},
  {11, 12.2, 12.3},
  {11.3, 11.9, 12.5},
  {13.1, 12.1, 12.9},
  {13.7, 13.4, 14.1},
  {14.6, 15.6, 16.2},
  {15.9, 16.6, 17.4},
  {15.4, 17.4, 18.9},
  {14.8, 17.6, 18.9},
  {15.3, 18, 17.2},
  {15.6, 17.6, 18.7},
  {15.9, 17.5, 18.6},
  {15, 16.6, 17.4},
  {11.8, 14.1, 15},
  {10.7, 13.2, 13.6},
  {11.2, 13.3, 12.6},
  {11.4, 13, 12.5},
  {11.7, 12.9, 12.5},
  {11.9, 12.2, 12.6},
  {10.7, 11.7, 12.5},
  {10.1, 11.5, 11.4},
  {9.4, 11.4, 10.5},
  {10, 11, 10},
  {9.2, 10.6, 9.7},
  {9, 10.3, 10.6},
  {9.4, 10.4, 10.8},
  {10.6, 10.7, 11},
  {14, 12.9, 11.4},
  {15, 15.1, 13.5},
  {16, 17, 17.9},
  {17.6, 17.5, 20.6},
  {18.7, 19.3, 22.4},
  {19.6, 20.7, 23.6},
  {19.6, 21.5, 22.9},
  {19.4, 21.2, 22.6},
  {18.7, 21.1, 21.2},
  {16.4, 19.5, 19},
  {14.4, 17.6, 16.5},
  {13, 16.5, 14.5},
  {12.3, 15.5, 13.8},
  {12, 15.3, 13.1},
  {12.9, 15.4, 12.6},
  {12.9, 15.3, 12.8},
  {13.7, 14.7, 13.1},
  {13.6, 14.3, 13.2},
  {12.6, 13.4, 12.7},
  {11.6, 13, 11.9},
  {11.8, 12.9, 11.2},
  {11.3, 12.8, 10.6},
  {11.7, 12.8, 10.5},
  {13, 13.1, 11},
  {16.1, 14.3, 13.8},
  {17.5, 16.9, 17.3},
  {17.9, 18.1, 20.5},
  {19.5, 19.3, 22.8},
  {19.9, 20.9, 24.5},
  {20.6, 22.3, 24.6},
  {20.7, 22.8, 24.1},
  {19.6, 22.6, 23.8},
  {18.6, 21.5, 22.6},
  {17.4, 20.7, 21.2},
  {16.9, 18.3, 18.7},
  {15.6, 17.2, 16.7},
  {14, 16.1, 15.4},
  {13.5, 15.6, 14.4},
  {13.4, 15.1, 13.9},
  {13.3, 15.1, 13.7},
  {13, 14.9, 13.1},
  {13, 14.3, 12.6},
  {12.5, 14.3, 12.3},
  {12.6, 14, 12.1},
  {12.1, 13.6, 11.7},
  {11.8, 13, 11.6},
  {12, 13.3, 12.5},
  {13.6, 13.6, 13.1},
  {17.7, 15.1, 13.7},
  {18.7, 17.3, 16.7},
  {18.8, 18.8, 20.9},
  {19.9, 19.9, 23.5},
  {20.8, 21.6, 25.3},
  {21.3, 22.8, 25.5},
  {21.4, 23.5, 24.2},
  {20.7, 23, 23.8},
  {19.8, 22.1, 23.2},
  {17.8, 20.5, 21.3},
  {17.1, 18.6, 19.9},
  {16.9, 17.8, 18.2},
  {16.9, 17.5, 17.3},
  {16.3, 17.8, 17.1},
  {15.9, 17.5, 16.9},
  {15.7, 17.1, 17},
  {15.4, 16.9, 16.8},
  {16, 16.6, 16.7},
  {15.7, 16.4, 16.4},
  {15.4, 16.3, 16.2},
  {15.4, 16, 16.1},
  {15.1, 15.9, 15.9},
  {14.6, 15.8, 16},
  {15.3, 15.9, 16.4},
  {17, 16.5, 17.7},
  {16.9, 17.2, 19.1},
  {18.1, 18.1, 20.3},
  {18.5, 19.1, 21.4},
  {18.1, 19.4, 21.3},
  {17.3, 19.3, 21},
  {17.1, 19.1, 21.5},
  {17, 19.2, 21.6},
  {16.5, 18.8, 21},
  {16.4, 18.2, 20.1},
  {16, 17.4, 19},
  {14.2, 17, 17.6},
  {14.8, 16.9, 16.4},
  {14.1, 16.3, 15.3},
  {15.1, 16.1, 14.6},
  {14.6, 16, 14.1},
  {14.2, 16.4, 13.5},
  {13.1, 16.2, 12.9},
  {12.5, 16.1, 13},
  {12.1, 15.9, 13.3},
  {12.8, 15.3, 12.9},
  {12.8, 14.8, 13.3},
  {13.4, 14, 13.7},
  {13.9, 13.4, 14.3},
  {14, 13.7, 15.7},
  {13.6, 14.5, 17.6},
  {13.5, 16.1, 18.2},
  {13, 14.1, 16.9},
  {12.7, 13.2, 16},
  {12.1, 12.7, 15.4},
  {11.6, 11.9, 14.7},
  {11.3, 11.4, 14.4},
  {10.6, 11, 14},
  {10.1, 10.5, 13.4},
  {9.6, 10, 12.8},
  {9.1, 9.6, 12.2},
  {8.7, 9, 11.9},
  {8.3, 8.7, 12},
  {7.9, 8.3, 11.8},
  {7.5, 8, 10.8},
  {7, 7.9, 10.2},
  {6.8, 7.8, 10},
  {6.6, 7.5, 9.9},
  {6.5, 7.5, 9.6},
  {6.5, 7.4, 9.5},
  {6.4, 7.3, 9.4},
  {6.5, 7.3, 9.5},
  {6.6, 7.4, 9.6},
  {7, 7.6, 9.8},
  {7.3, 7.8, 10.3},
  {8.1, 8.5, 11.5},
  {8.4, 9.9, 12.3},
  {8.6, 10.9, 13.1},
  {9.6, 10.9, 14.3},
  {10.4, 11.3, 16.1},
  {10.7, 11.6, 16.3},
  {10.9, 12.1, 15.3},
  {10.4, 10.6, 13.6},
  {9.5, 10.1, 13.2},
  {9.1, 10, 12.6},
  {9, 10.2, 12.1},
  {8.9, 10.3, 11.7},
  {8.7, 10.1, 11.4},
  {8.6, 9.7, 11.2},
  {8.5, 9.5, 11},
  {8.4, 9.2, 10.9},
  {8.2, 9, 10.7},
  {7.9, 8.9, 10.6},
  {7.8, 8.7, 10.4},
  {7.8, 8.7, 10.4},
  {8.1, 8.8, 10.4},
  {8.8, 9.6, 10.8},
  {9.3, 10.3, 11.3},
  {9.7, 11, 12.3},
  {10.1, 11.4, 13.9},
  {10.8, 12.3, 15.2},
  {11, 12.9, 16.6},
  {11.2, 13.4, 16.5},
  {11.8, 13.5, 17.2},
  {11.7, 14.2, 17.3},
  {11.4, 13.9, 16.1},
  {11, 12.9, 15},
  {10.2, 12.3, 14.6},
  {9.4, 11.9, 13.9},
  {9.5, 11.6, 13.3},
  {9.8, 11.4, 13},
  {9.8, 11.2, 12.9},
  {9.8, 10.9, 12.8},
  {9.8, 10.9, 12.8},
  {9.7, 10.7, 12.6},
  {9.7, 10.6, 12.3},
  {9.6, 10.5, 12.1},
  {9.5, 10.4, 12},
  {9.6, 10.4, 11.8},
  {9.5, 10.4, 11.8},
  {9.9, 11.2, 12.2},
  {10.9, 12.3, 13.1},
  {11.6, 12.9, 15.1},
  {12.2, 14.8, 16.6},
  {13.5, 14.7, 18.4},
  {13.6, 14.9, 19.5},
  {14.9, 16.4, 19.9},
  {15.5, 17.3, 19.4},
  {14.4, 17.4, 18},
  {13, 16.9, 17.5},
  {12.2, 15.3, 16.7},
  {11.9, 13.4, 14.9},
  {11.7, 12.4, 13.5},
  {11.6, 12.1, 12.5},
  {11, 11.9, 11.8},
  {10.3, 11.9, 11.4},
  {10.3, 11.8, 11.1},
  {10, 11.8, 10.8},
  {9.5, 11.3, 10.7},
  {8.9, 10.4, 10.5},
  {8.4, 9.8, 9.8},
  {8.6, 10.1, 9.9},
  {9, 9.8, 10.2},
  {9.4, 10.2, 10.3},
  {10.3, 11.4, 11},
  {11.2, 11.9, 12.6},
  {12.5, 13, 15.7},
  {13.7, 14.9, 18.4},
  {13.9, 15.2, 19.1},
  {14.9, 17.1, 19.1},
  {15.6, 17.7, 18.4},
  {14.8, 17.4, 17.8},
  {14.4, 17, 17.2},
  {14.5, 17, 16.9},
  {13.1, 15.1, 16.3},
  {12.2, 14.2, 15.2},
  {11.7, 13.3, 14.3},
  {11.8, 13.1, 13.8},
  {11.4, 13.1, 13.5},
  {11.6, 12.7, 13.1},
  {11.5, 12.8, 13.3},
  {11, 13.1, 13.2},
  {10.8, 12.8, 13.2},
  {10.6, 12.5, 13},
  {10.5, 12.2, 13},
  {10, 11.9, 12.7},
  {9.9, 11.6, 12.6},
  {9.8, 11.7, 12.5},
  {10.7, 12.4, 12.7},
  {11.2, 12.5, 13.2},
  {12.3, 13.6, 13.9},
  {12.7, 14.6, 15.7},
  {13.4, 15.9, 18.6},
  {14, 16.9, 18.8},
  {14.1, 17.6, 18.9},
  {14.5, 17.4, 20.2},
  {15.2, 17.5, 19.2},
  {15.3, 17, 17.9},
  {13.4, 16.1, 16.5},
  {11.2, 14.2, 14.4},
  {10.3, 13.3, 12.6},
  {10, 12.2, 11.6},
  {10.3, 12.2, 10.9},
  {10.4, 11.8, 10.3},
  {9.3, 11.1, 9.8},
  {9.8, 11.4, 9.4},
  {9.7, 11.8, 9.2},
  {10.3, 11.8, 9.4},
  {10.5, 11.7, 9.4},
  {9, 11.4, 9.2},
  {8.6, 11.1, 9.2},
  {8.9, 10.5, 9.7},
  {10.6, 10.7, 9.9},
  {12.1, 12, 11.1},
  {13.6, 14.9, 13.8},
  {15.4, 15.3, 17.4},
  {15.8, 16.8, 19.9},
  {16.6, 18.4, 20.7},
  {17, 19.3, 20.3},
  {16.5, 19.4, 19.9},
  {15.9, 18.9, 20.1},
  {14.9, 18.2, 19.3},
  {13.4, 16, 18},
  {12.8, 14.5, 16.7},
  {11.6, 14, 15.6},
  {12.3, 13.5, 15.2},
  {11.1, 13.4, 14.9},
  {10.6, 12.7, 14.6},
  {10, 12.4, 14.4},
  {10.2, 12.3, 13.8},
  {10.8, 11.8, 13.8},
  {10.6, 11.4, 13.7},
  {9.9, 12.1, 12.9},
  {9.5, 12.4, 12.8},
  {9.7, 11.9, 12.2},
  {10.1, 11.3, 11.3},
  {10.7, 11.7, 11.2},
  {14.1, 12.8, 13},
  {15.7, 15.1, 16.8},
  {15.8, 17.3, 19.3},
  {17.1, 17.8, 21.6},
  {17.8, 19.3, 22.5},
  {18.4, 20.7, 22.4},
  {18.6, 21.4, 21.5},
  {18.2, 20.9, 21},
  {17.1, 19.4, 19.6},
  {15.4, 17.2, 18.3},
  {13.1, 16.1, 16},
  {12.5, 15.3, 14.3},
  {11.6, 14.7, 13.4},
  {11.1, 13.7, 12.6},
  {11, 13.1, 11.8},
  {10.4, 13.1, 11.2},
  {10.3, 12.1, 10.9},
  {9.6, 11.1, 10.9},
  {9.5, 11.4, 10.7},
  {9.6, 10.7, 10.5},
  {9.7, 10.5, 9.6},
  {9.1, 10.4, 9},
  {9.4, 10.3, 8.6},
  {10.7, 10.9, 9.4},
  {14.1, 12.5, 11.3},
  {15.5, 14.2, 14.3},
  {15.9, 15.9, 17.8},
  {16.7, 17.1, 20},
  {17.3, 18.4, 20.5},
  {17.1, 18.5, 20.6},
  {17.6, 19.7, 21.4},
  {17, 19, 19.3},
  {14.7, 16.6, 18.4},
  {14.2, 16.2, 17.1},
  {13.3, 14.8, 16.1},
  {12.5, 13.6, 15.2},
  {11.6, 13.1, 13.5},
  {11.4, 12.4, 12.2},
  {10.5, 12.1, 11.1},
  {10.1, 11.9, 10.4},
  {10.7, 11.3, 9.6},
  {9.8, 11.2, 9},
  {9.4, 10.8, 8.4},
  {9.6, 10.6, 8.2},
  {9.2, 10.6, 7.9},
  {9.2, 10.4, 8.2},
  {9.3, 10.4, 9.2},
  {9.9, 10.6, 9.4},
  {13.3, 11.6, 9.9},
  {15.1, 14.8, 12.5},
  {15.7, 16.4, 16.4},
  {17.2, 17.3, 19.8},
  {17.8, 18.8, 21.3},
  {18.3, 20.3, 22.5},
  {18.7, 20.5, 21.4},
  {16.9, 20, 20.6},
  {16.1, 19, 20.3},
  {14.7, 17.3, 18.2},
  {13.9, 16, 16},
  {12, 15.2, 14},
  {11.7, 14.3, 12.9},
  {11.4, 13.7, 12.2},
  {11.5, 13.5, 11.8},
  {12.4, 14, 12.4},
  {12.1, 14.2, 12.5},
  {11.1, 14.1, 12.5},
  {11.2, 13.7, 12.7},
  {11.4, 12.9, 12.8},
  {11.3, 12.5, 12.4},
  {11.2, 12.7, 12.2},
  {11.4, 13, 12},
  {12.2, 13.2, 12.4},
  {13.2, 13.6, 13.4},
  {14.3, 14.2, 14.7},
  {14.6, 14.5, 16.2},
  {15.1, 15.3, 17.8},
  {15.6, 16.2, 19},
  {15.5, 16.8, 19.3},
  {15.3, 16, 19.5},
  {15.2, 15.3, 19.2},
  {14.3, 14.4, 18.7},
  {13.7, 14.1, 18},
  {12.7, 13.7, 16.6},
  {12.4, 13.5, 15.6},
  {12.6, 13.4, 15},
  {12.5, 13.2, 14.6},
  {12.1, 13, 14.3},
  {11.4, 12.7, 13.9},
  {11.2, 12.5, 13.2},
  {10.6, 12.4, 12.4},
  {10.4, 12, 12.1},
  {11.5, 12.1, 12.1},
  {11.6, 12.5, 12.3},
  {11.4, 11.9, 12.1},
  {11.2, 11.4, 11.9},
  {11.8, 11.8, 11.9},
  {13.7, 12.7, 12.7},
  {14.7, 14.9, 14.9},
  {15.7, 15.4, 18.9},
  {16.5, 16.8, 20.6},
  {17.4, 18.5, 21.9},
  {18.4, 19.8, 21.8},
  {18.2, 20.2, 20.4},
  {16.4, 19.2, 19.8},
  {15, 17.9, 18.9},
  {15, 16.5, 18.3},
  {14.9, 16, 17.4},
  {14.5, 16, 16.8},
  {13.8, 15.8, 15.8},
  {14.1, 15.5, 15},
  {13.9, 15.8, 14.3},
  {12.9, 15.5, 13.8},
  {13.7, 15.5, 13.7},
  {13.8, 15.4, 13.7},
  {13.6, 15.1, 13.7},
  {13.5, 15.3, 13.6},
  {13.2, 14.2, 13.7},
  {13.4, 14, 13.7},
  {13.3, 13.9, 13.6},
  {13.1, 13.8, 13.8},
  {13.2, 13.8, 14},
  {14.2, 13.8, 14.4},
  {13.6, 14.7, 14.9},
  {14.1, 15, 15.8},
  {13.5, 15.1, 16.6},
  {13.6, 13.6, 17},
  {13.6, 12.5, 17.5},
  {13.7, 12, 16.9},
  {12.7, 13.2, 14.4},
  {12.1, 12.4, 14.1},
  {10.6, 10.9, 12.4},
  {9.4, 10.7, 11},
  {9.3, 11.2, 10.8},
  {8.9, 11.5, 10.4},
  {8.4, 10.7, 10},
  {7.8, 9.9, 9.9},
  {7.7, 9.7, 10.2},
  {7.6, 9.3, 10.4},
  {8.1, 8.6, 10.3},
  {7.2, 7.8, 10.1},
  {6.3, 8.7, 9.9},
  {6, 8.1, 9.7},
  {6.4, 7.6, 9.4},
  {6.6, 7.4, 9.4},
  {10.3, 8.5, 10.5},
  {11.9, 10.8, 12.4},
  {13.2, 13, 15.2},
  {13.6, 14.5, 17.5},
  {14.6, 15.4, 18.2},
  {15.2, 16.1, 18.9},
  {15.8, 16.6, 19.5},
  {15.3, 16.6, 19.7},
  {14.3, 16.1, 17},
  {9.4, 13.3, 13.2},
  {7.9, 11.3, 10.1},
  {8.4, 10.7, 8.8},
  {8.1, 9.9, 8.7},
  {8.9, 9, 8.5},
  {9.7, 8.7, 7.9},
  {8.9, 8.7, 8.3},
  {8.6, 8.8, 8.4},
  {8.6, 8.2, 8.8},
  {8.6, 8.3, 8.9},
  {8.4, 7.9, 9.1},
  {8.1, 7.3, 9.1},
  {7.8, 7.3, 9.1},
  {8, 7.2, 9},
  {8.9, 7.7, 9.3},
  {9.7, 8, 10.9},
  {11.4, 11.1, 13},
  {11.8, 12.9, 15.4},
  {12.4, 13.7, 17.1},
  {13, 14.7, 17.2},
  {13.4, 15.6, 15.9},
  {13.4, 15.6, 17.4},
  {12.7, 16.1, 16.6},
  {11.7, 15.1, 15.6},
  {10.5, 12.9, 13.7},
  {10.2, 11.9, 12.1},
  {10.4, 11.5, 11.1},
  {10.1, 10.7, 10.4},
  {10.2, 10.1, 10.2},
  {9.4, 10.1, 10.1},
  {9.3, 10.2, 10.1},
  {9.3, 9.9, 10.1},
  {8.8, 9.6, 10},
  {8.9, 9.5, 9.9},
  {8.8, 9.4, 10},
  {8.6, 9.4, 10.1},
  {8.5, 9.4, 10.2},
  {8.4, 9.4, 10.1},
  {8.6, 9.7, 10.4},
  {9, 9.9, 10.6},
  {9, 10, 10.9},
  {8.9, 10.3, 11.2},
  {8.8, 10.3, 11.2},
  {8.8, 10.1, 11.2},
  {9, 10.1, 11.1},
  {8.8, 10, 11.4},
  {8.6, 9.8, 11.5},
  {8.7, 8.8, 11.4},
  {8.6, 8.1, 10.7},
  {8.4, 7.9, 10.3},
  {7.9, 7.6, 10.2},
  {7.5, 7.3, 9.9},
  {6.6, 7.3, 8.9},
  {5.9, 7.2, 8.3},
  {6.3, 7, 7.9},
  {6.1, 6.8, 7.5},
  {5.9, 6.3, 7.6},
  {5.7, 6, 7.6},
  {5.6, 5.8, 7.6},
  {5.4, 5.9, 7.6},
  {5.3, 5.9, 7.5},
  {5.5, 6.1, 7.6},
  {5.5, 6.4, 7.7},
  {5.8, 6.8, 8.1},
  {7.2, 7.4, 8.6},
  {6.7, 7.3, 8.8},
  {6.9, 7.5, 8.8},
  {7.3, 7.3, 9.2},
  {7.2, 7.1, 9.4},
  {7.1, 7.2, 9.6},
  {6.7, 7.5, 9.6},
  {7.1, 7.6, 9.4},
  {7.9, 7.6, 9.4},
  {7.8, 7.6, 9.2},
  {7.4, 7.6, 9},
  {6.8, 7.5, 9},
  {6.4, 7.6, 9.1},
  {6.9, 7.7, 9.1},
  {7.6, 7.7, 8.8},
  {7.6, 7.7, 8.3},
  {7.7, 7.5, 7.8},
  {7.6, 7, 8.1},
  {7.6, 6.8, 8.2},
  {7.4, 6.9, 8.1},
  {6.5, 6.7, 8.1},
  {6.2, 7, 7.5},
  {6.9, 7.6, 7.8},
  {8.3, 8.2, 8.2},
  {8.7, 8.5, 9.6},
  {8.8, 9, 10},
  {9.4, 9.1, 10.9},
  {9, 9.4, 11.4},
  {8.9, 9.3, 11.6},
  {9.8, 8.9, 12},
  {9.2, 9.2, 11.6},
  {8.5, 8.9, 11.3},
  {8, 8.4, 10.3},
  {7.5, 8.2, 9.8},
  {7.2, 8.3, 9.7},
  {6.9, 8.3, 9.4},
  {5.7, 7.9, 8.4},
  {5.4, 7.6, 7.6},
  {5.7, 7.6, 7.5},
  {5.3, 7.4, 7.5},
  {5, 7.4, 7.3},
  {4.7, 7.5, 7.3},
  {5.2, 7.7, 7.3},
  {5.3, 7.5, 7.2},
  {5.4, 7.5, 7.1},
  {6.3, 7.5, 7.2},
  {6.9, 7.6, 7.3},
  {6.9, 7.9, 7.7},
  {7, 8.5, 8.3},
  {7.4, 9.3, 9},
  {7.1, 10.1, 9.5},
  {7.8, 10.5, 10},
  {8.9, 10.5, 11.1},
  {9, 10.5, 11.3},
  {8.9, 10.1, 11.1},
  {8.8, 9.9, 10.9},
  {8.8, 9.6, 10.7},
  {8.7, 9.2, 10.5},
  {8.7, 9.2, 10.4},
  {8.8, 9.3, 10.4},
  {8.7, 9.4, 10.4},
  {8.4, 9.3, 10.3},
  {8.4, 9.3, 10.2},
  {8.8, 9.7, 9.9},
  {8.3, 9.4, 9.9},
  {8.4, 9.5, 10},
  {8.3, 9.4, 10.1},
  {8.3, 9.5, 10.1},
  {8.5, 9.5, 10.2},
  {8.7, 9.6, 10.1},
  {9, 9.8, 10.1},
  {9.8, 10.3, 10.6},
  {10.2, 11.1, 11},
  {10.2, 11.5, 11.3},
  {11.3, 11.2, 11.6},
  {11.8, 11.5, 12},
  {11.7, 11.9, 12.2},
  {12, 11.8, 12.3},
  {10.8, 11.6, 12.1},
  {10.6, 11.4, 12},
  {10.5, 10.9, 11.8},
  {10.4, 10.5, 11.6},
  {10, 10.1, 11.2},
  {10.4, 10.1, 11.2},
  {10.5, 10.3, 11.1},
  {10.5, 10.2, 11},
  {10.2, 10.3, 10.9},
  {9.5, 10.2, 10.9},
  {9.5, 10, 10.9},
  {9.5, 9.9, 10.9},
  {9.7, 9.7, 10.9},
  {9.6, 10, 10.8},
  {9.3, 10, 10.9},
  {9.2, 10, 11},
  {9.3, 10.1, 11.1},
  {9.7, 10.5, 11.5},
  {9.9, 10.8, 11.9},
  {10.3, 11.4, 12.1},
  {10, 11.4, 12.3},
  {10, 12.1, 12.4},
  {10.6, 12.4, 12.5},
  {10.8, 12.3, 12.6},
  {10.4, 12.2, 12.6},
  {10, 11.6, 12.6},
  {9.4, 11.1, 12.3},
  {9.1, 10.6, 11.9},
  {8.8, 10.4, 11.8},
  {9.1, 10.2, 11.6},
  {9.4, 10.1, 11.6},
  {9.2, 10.1, 11.5},
  {8.8, 9.9, 11.2},
  {8, 9.5, 10.5},
  {9, 9.6, 10.6},
  {8.8, 9.8, 10.6},
  {9.2, 9.8, 10.5},
  {8.4, 9.9, 10.4},
  {8.8, 10, 10.4},
  {8.5, 9.9, 10.4},
  {8.7, 9.9, 10.5},
  {9.1, 10, 10.8},
  {9.4, 10.7, 11.3},
  {10.2, 12.3, 11.9},
  {11.7, 14.1, 13.8},
  {12.9, 13.9, 16.3},
  {12.2, 14, 16.7},
  {12.5, 14.4, 16.8},
  {12.6, 14.3, 16.6},
  {12.1, 13.5, 16.2},
  {11.5, 12.2, 14.9},
  {10.9, 11.5, 13.5},
  {10.7, 11.5, 12.9},
  {10.7, 11.3, 12.3},
  {10.4, 11.3, 12},
  {10.3, 11.1, 11.9},
  {10.2, 11.1, 11.7},
  {10.2, 10.9, 11.5},
  {9.9, 11, 11.4},
  {9.7, 11.1, 11.5},
  {9.8, 11.1, 11.5},
  {9.8, 11.1, 11.6},
  {9.7, 10.9, 11.6},
  {9.6, 10.9, 11.6},
  {9.3, 10.5, 11.8},
  {10.5, 10.5, 12},
  {11.8, 12, 14.2},
  {12.5, 14.1, 16.7},
  {12.1, 14.7, 18.4},
  {13.4, 15.8, 19.3},
  {14.4, 16.8, 19.4},
  {14.5, 17.7, 18.4},
  {13.4, 16.7, 17},
  {11.9, 15.2, 16.4},
  {10.8, 13.4, 14.6},
  {9.3, 11.8, 12.7},
  {9.4, 11.7, 11.6},
  {9.3, 11.2, 11.8},
  {9.2, 10.9, 11.9},
  {9, 11.1, 11.7},
  {9.8, 10.8, 11},
  {9.4, 10, 10.5},
  {9.7, 10.5, 11},
  {9.7, 10.6, 11.2},
  {8.7, 10.8, 11},
  {7.7, 10.8, 11.2},
  {8.9, 10.7, 11.4},
  {8.8, 10.5, 11.6},
  {9.5, 11, 11.8},
  {9.9, 11.5, 12.3},
  {10.3, 11.7, 12.8},
  {10.9, 12.2, 13.7},
  {11.7, 12.7, 15.1},
  {12.7, 13.9, 16.5},
  {12.8, 14.6, 17.2},
  {13.6, 15.8, 17.7},
  {13.2, 15.8, 15.8},
  {12.2, 14.9, 15.3},
  {8.7, 12.6, 13.5},
  {7.8, 11.8, 11.3},
  {7.9, 11.3, 9.9},
  {8.4, 11.2, 9.3},
  {8.2, 10.9, 8.6},
  {7.8, 10.4, 8.8},
  {7.4, 9.6, 9},
  {7.7, 10.3, 8.8},
  {8.1, 9.8, 9.1},
  {7.5, 9.1, 9},
  {7.4, 8.9, 8.7},
  {7, 8.1, 8.2},
  {6.7, 7.3, 7.3},
  {6.5, 7.3, 6.9},
  {7.9, 7.4, 7.3},
  {10.3, 8.4, 8.8},
  {12, 9.7, 12.2},
  {13, 12.5, 15.7},
  {13.9, 14.1, 16.5},
  {12.2, 15, 17.7},
  {13, 15.7, 18.7},
  {13.9, 16.1, 18.3},
  {13.1, 16.1, 17.4},
  {11.2, 14.6, 15.4},
  {9.6, 11.8, 12.5},
  {7.5, 10.4, 10.3},
  {7, 9.7, 9},
  {6.7, 10, 8.8},
  {6.6, 9.5, 8.1},
  {6.6, 9.3, 7.3},
  {6.7, 8.3, 6.6},
  {6.6, 7.8, 6.1},
  {6.1, 7.2, 5.5},
  {6.8, 6.4, 4.9},
  {6, 5.6, 4.4},
  {5.6, 5.6, 3.8},
  {5.5, 5.4, 3.5},
  {4.9, 5.6, 3.1},
  {5.8, 6.1, 3.6},
  {8.3, 6.8, 5.4},
  {10.5, 8.3, 7.8},
  {10.7, 10.3, 11},
  {11.5, 11.8, 14.6},
  {12.3, 13, 16.6},
  {12.5, 14.4, 16.4},
  {12.3, 14.8, 15.7},
  {10.3, 14, 15},
  {9.1, 12.7, 13.3},
  {8.3, 10.4, 12.2},
  {8.5, 9.2, 10.4},
  {8.2, 8.4, 9},
  {8.7, 8, 8},
  {8.5, 7.7, 8.2},
  {8, 8.4, 8.5},
  {7.9, 8.5, 8.8},
  {7.4, 8.1, 8.8},
  {6.1, 8, 8.7},
  {5.9, 8.1, 8.4},
  {5.2, 7.9, 7.8},
  {4.7, 7.2, 7.2},
  {4.1, 6.8, 6.9},
  {4.1, 6.6, 6.2},
  {4.8, 6.6, 5.7},
  {7.7, 7.1, 6.6},
  {9.6, 8.3, 8.7},
  {10.7, 10.5, 12},
  {11.2, 12, 14.6},
  {12, 13.3, 15.9},
  {12.6, 14.4, 16.5},
  {12.8, 14.6, 16},
  {11.3, 14.1, 15},
  {9.8, 13, 13.7},
  {8.5, 10.9, 11.5},
  {8.7, 9.5, 9},
  {8.1, 8.1, 7.6},
  {7, 7.4, 7},
  {5.8, 7.6, 6},
  {5.1, 7.1, 5.5},
  {4.8, 6.6, 5},
  {4.7, 6.7, 4.5},
  {4.9, 6.5, 4.2},
  {4.6, 6.8, 3.8},
  {4.1, 6.3, 4.1},
  {4.2, 6, 5.2},
  {4.3, 5.7, 5.7},
  {4.3, 5.8, 5.6},
  {4.4, 5.7, 5.3},
  {7.1, 6.7, 5.4},
  {10.1, 8.2, 5.7},
  {11.3, 10.8, 7.7},
  {12.5, 11.2, 11.7},
  {13.2, 13, 15.5},
  {13.8, 14.5, 17.7},
  {14.3, 15.7, 18.2},
  {13.7, 15.3, 16.8},
  {12, 14.1, 15.2},
  {8.3, 11.4, 12.3},
  {7.3, 10.4, 9.5},
  {6.3, 9.9, 8.1},
  {6.1, 9.1, 7.2},
  {6.2, 8.3, 6.4},
  {6.2, 7.9, 5.8},
  {5.8, 7.8, 5.5},
  {5.7, 7.7, 4.7},
  {5.4, 7.3, 4.4},
  {5.6, 7.1, 4.7},
  {5.2, 7.2, 5.5},
  {4.9, 6.7, 6},
  {5, 6.4, 5.9},
  {4.8, 6.1, 5.7},
  {5.3, 6, 5.6},
  {7.7, 6.8, 5.5},
  {10.7, 7.9, 6.1},
  {12.4, 11.1, 8.1},
  {13.6, 12.3, 12.3},
  {14, 13.5, 16.2},
  {14.5, 15.2, 18.4},
  {14.8, 15.8, 18.8},
  {14.4, 16, 17.5},
  {12, 15.2, 15.7},
  {9.2, 12.1, 13.1},
  {8.1, 10.3, 10.6},
  {7.2, 9.8, 9},
  {6.5, 8.8, 8},
  {6.6, 8.5, 6.9},
  {6.6, 8.4, 6.3},
  {7.4, 8.3, 5.8},
  {7.2, 8.4, 5.2},
  {7.1, 8.2, 4.9},
  {6, 7.9, 4.8},
  {5.7, 7.4, 5.4},
  {5.6, 7.1, 6.2},
  {5.3, 6.7, 6.3},
  {5.1, 6.4, 6.1},
  {6, 6.4, 5.8},
  {9, 7.6, 5.8},
  {12.4, 9.3, 6.3},
  {13.3, 11.4, 8.3},
  {14.8, 12, 13},
  {15, 14.2, 17.1},
  {15.6, 15.5, 19.1},
  {15.6, 16.4, 19.8},
  {14.9, 16.6, 18.1},
  {13.4, 16, 15.8},
  {9.5, 12.1, 12.5},
  {8.5, 10.8, 10.3},
  {7.9, 10.4, 8.8},
  {7.8, 10.8, 7.8},
  {8.3, 10.1, 7},
  {8.6, 9.3, 6.5},
  {8.8, 8.7, 6},
  {8.7, 8.4, 5.6},
  {7.8, 8.2, 5.1},
  {6.4, 7.7, 5},
  {6.6, 7.3, 4.8},
  {7.1, 7, 4.8},
  {8.2, 6.8, 5.5},
  {8.1, 6.4, 5.6},
  {8.4, 7.2, 6.1},
  {8.5, 8.3, 6.6},
  {8.3, 9.1, 7.5},
  {8, 10.5, 8.5},
  {7.8, 11.7, 10},
  {7.7, 12.2, 11.8},
  {8.3, 12.2, 12.1},
  {8.7, 11.9, 12},
  {8.4, 11.4, 11.7},
  {8.2, 10.2, 11.5},
  {7.8, 9, 11.3},
  {7.6, 8.9, 10.9},
  {7.6, 9.6, 10.5},
  {7.5, 9.6, 10.2},
  {7.4, 9.6, 10},
  {7.3, 8.9, 9.9},
  {7, 9, 9.7},
  {6.9, 8.9, 9.6},
  {6.8, 8.5, 9.6},
  {6.6, 8.5, 9.5},
  {6.4, 8.2, 9.4},
  {6.1, 8.2, 9.1},
  {5.7, 8, 9.4},
  {5.8, 8, 9.5},
  {5.9, 8, 9.4},
  {6.1, 8, 9.7},
  {6, 8.3, 9.8},
  {6.1, 9.1, 9.9},
  {6, 9.9, 10.1},
  {6.1, 10.7, 10.4},
  {6.4, 11.3, 10.9},
  {7.8, 11.8, 11.1},
  {7.9, 11.1, 10.9},
  {7.8, 9.6, 10.8},
  {5.1, 8.2, 10.4},
  {3.7, 7.1, 8.8},
  {3.7, 6.7, 6.9},
  {3.4, 6.4, 5.7},
  {3.4, 6.9, 5.1},
  {3.3, 6.9, 4.3},
  {3.2, 7.1, 3.7},
  {3.1, 7, 3.3},
  {3.5, 6.9, 2.8},
  {3.7, 6.8, 3.5},
  {4.1, 6.8, 4.2},
  {4.8, 6.8, 4.4},
  {4.7, 6.7, 4.1},
  {3.8, 6.6, 3.7},
  {4.9, 6.9, 4.2},
  {7, 7.4, 5.4},
  {7.9, 8, 6.6},
  {8.1, 8.9, 8.2},
  {7.8, 9.7, 10.3},
  {7.7, 10.1, 12.2},
  {7.1, 10, 11.4},
  {7.9, 9.5, 11.2},
  {7.5, 9.7, 11.4},
  {7, 9.4, 11.1},
  {6.4, 8.6, 10},
  {6.2, 8.3, 9.7},
  {6.3, 8.2, 9.5},
  {6.4, 8.1, 9.2},
  {6.4, 8, 8.9},
  {6.4, 7.9, 8.8},
  {6.5, 7.7, 8.4},
  {6.5, 7.5, 8.3},
  {6.5, 7.3, 8.3},
  {6.7, 7.2, 8},
  {6.6, 7, 7.9},
  {6.5, 7.3, 7.9},
  {6.3, 7.4, 7.8},
  {6.3, 7.4, 7.6},
  {6.4, 7.4, 8},
  {6.7, 7.6, 8.3},
  {7.1, 7.6, 8.7},
  {7.1, 8.1, 9.3},
  {7.5, 8.3, 9.7},
  {7.8, 8.3, 9.9},
  {8.1, 8.6, 10},
  {8, 8.7, 10.2},
  {7.8, 8.7, 10.3},
  {7.8, 9, 10.3},
  {7.6, 8.6, 10.1},
  {7.7, 8.5, 10},
  {7.8, 8.5, 9.7},
  {7.7, 8.5, 9.7},
  {7.9, 8.3, 9.6},
  {8.1, 8.4, 9.7},
  {8.1, 8.4, 9.6},
  {8.2, 8.3, 9.6},
  {8.1, 8.3, 9.5},
  {8.1, 8.3, 9.5},
  {8.1, 8.2, 9.4},
  {8.1, 8.1, 9.4},
  {8, 8.2, 9.4},
  {8.1, 8.2, 9.4},
  {8.6, 8.4, 9.4},
  {9.3, 8.9, 9.9},
  {9, 9.3, 10.3},
  {9.3, 9.9, 11.2},
  {9.5, 10.3, 12.6},
  {10.6, 10.8, 13.6},
  {12, 11.7, 15},
  {12.5, 12.2, 16.2},
  {11.5, 13, 15.2},
  {10.1, 12, 13},
  {8.3, 10.9, 12.1},
  {8.1, 10.7, 11.6},
  {8.3, 10.8, 11.5},
  {8.8, 10.8, 11.4},
  {9, 10.6, 10.9},
  {9, 10.1, 10.4},
  {9, 9.5, 10.5},
  {8.3, 8.3, 10.1},
  {6.7, 9.1, 10.3},
  {6.7, 8.9, 10.1},
  {6.3, 8, 9.5},
  {5.9, 7.9, 9.5},
  {5.9, 7.2, 9.2},
  {6.5, 7.4, 9.2},
  {7.5, 7.6, 9.2},
  {8.5, 9, 9.5},
  {9.5, 10, 9.8},
  {10.7, 11.5, 11.1},
  {11.4, 11.8, 12.2},
  {11.7, 12.8, 14.7},
  {11.8, 13.6, 16.3},
  {12.5, 14.1, 17.2},
  {11.8, 15, 16.2},
  {11.1, 13.6, 14.3},
  {10.1, 11.5, 12.1},
  {9.9, 11, 10.6},
  {9.8, 10.2, 10.5},
  {9.6, 10.5, 10.4},
  {9.3, 10.4, 10.4},
  {9.6, 10.7, 10.4},
  {9.8, 11, 10.3},
  {9.7, 10.7, 10.3},
  {9.7, 10.2, 10.3},
  {9.7, 10.3, 10.3},
  {9.6, 10.2, 10.3},
  {9.6, 10.3, 10.3},
  {9.7, 10.3, 10.3},
  {9.7, 10.1, 10.4},
  {9.8, 10.2, 10.5},
  {10, 10.3, 10.9},
  {10.1, 10.4, 11.5},
  {10.3, 10.8, 12.2},
  {11.4, 11.1, 13.3},
  {11.1, 11.7, 14.1},
  {11.5, 12.1, 14.7},
  {11.9, 12.6, 15},
  {12.2, 13.1, 14.9},
  {12.3, 13, 14.5},
  {12.1, 12.6, 13.7},
  {11.2, 12, 13.5},
  {10.7, 11.9, 13.4},
  {10.7, 11.9, 13.3},
  {10.7, 11.8, 13.2},
  {10.6, 11.7, 13.1},
  {10.6, 10.8, 12.5},
  {10.1, 10.6, 12.2},
  {10.1, 10.3, 11.7},
  {9.3, 10.3, 11.8},
  {7.9, 10.8, 11.5},
  {8.1, 11, 10.9},
  {8.4, 10.9, 10.6},
  {8.4, 10.5, 10.2},
  {8.6, 10.8, 10.1},
  {9.8, 10.3, 10.2},
  {10.9, 10.8, 10.8},
  {11.2, 13.2, 12.8},
  {13.1, 13.7, 15.2},
  {14.1, 15.2, 17.3},
  {13.7, 16.1, 17.7},
  {13.8, 16.6, 17.1},
  {12.6, 16.1, 16.2},
  {12.3, 14.2, 14.9},
  {10.6, 12.4, 14.4},
  {9.3, 11.5, 14.1},
  {9.4, 11.2, 13.7},
  {9.7, 11.9, 13.5},
  {10.1, 12.1, 13.3},
  {9.2, 11.9, 13.2},
  {9, 12, 13},
  {9.6, 11.7, 12.9},
  {9.7, 11.5, 12.8},
  {9.6, 11.4, 12.2},
  {8.6, 11.1, 11.1},
  {8.2, 10.6, 10.7},
  {8.4, 9.9, 10.8},
  {9, 10.3, 11.1},
  {9.3, 10.4, 11.3},
  {9.6, 10.6, 11.7},
  {10.2, 10.9, 12.8},
  {11.2, 11.9, 13.9},
  {11.4, 13.2, 15},
  {12.7, 13.5, 15.8},
  {12.9, 13.9, 15.7},
  {12.1, 13.7, 15},
  {11.4, 13.8, 14.7},
  {10.6, 12.9, 14.5},
  {10.2, 12.6, 13.9},
  {10.1, 12.1, 13.4},
  {10.1, 11.7, 13.1},
  {10, 12.1, 12.7},
  {9.9, 12, 12.6},
  {9, 11.6, 12.3},
  {8.1, 11.5, 11.8},
  {7, 10.9, 11},
  {7, 10.8, 10.7},
  {6.7, 10.8, 10.8},
  {6.5, 10.3, 10.9},
  {6.3, 10.1, 10.7},
  {6.5, 10.1, 10.4},
  {6.1, 9.6, 9.9},
  {7.1, 9.4, 9.2},
  {9, 9.6, 9.3},
  {11.8, 10.2, 10.6},
  {12.8, 12.6, 12.9},
  {14, 13.4, 15.3},
  {14.5, 15, 17.8},
  {14.7, 16, 18.8},
  {14.9, 16.5, 18.6},
  {13.9, 15.8, 17.3},
  {11.6, 14.5, 15.7},
  {10, 12, 13.5},
  {10.6, 11.1, 11.7},
  {10.7, 10.7, 10.7},
  {10.6, 10.9, 10.7},
  {10.6, 10.8, 11},
  {10.4, 11.1, 10.9},
  {10.4, 10.8, 10.6},
  {10.2, 10.6, 10.3},
  {9.9, 10.6, 10.5},
  {9.9, 10.1, 10.6},
  {9.6, 9.2, 9.9},
  {8.8, 8.9, 8.8},
  {7.3, 8.7, 8},
  {6.9, 8.3, 8},
  {7.1, 8.4, 7.5},
  {8.6, 8.4, 8.2},
  {12, 9.5, 9.2},
  {13.1, 11.1, 10.6},
  {13.9, 12.9, 15.2},
  {14.8, 14.6, 17.2},
  {15, 15.8, 19.2},
  {15, 16.6, 19.2},
  {13.8, 16, 17.1},
  {11.4, 13.9, 15.3},
  {9, 12.2, 13.1},
  {8.7, 11.1, 11.2},
  {7.8, 10.6, 10.2},
  {7.5, 9.8, 9.2},
  {8.7, 9.8, 8.7},
  {9, 9.9, 9.5},
  {8.2, 9.6, 9.9},
  {8.4, 9.4, 10.2},
  {7.9, 9, 10.3},
  {7.3, 8.7, 10.3},
  {7, 8.5, 10.3},
  {6.8, 8.3, 10.1},
  {6.7, 8.1, 9.8},
  {7, 8, 9.5},
  {7.3, 8.3, 9.2},
  {9.3, 8.7, 9},
  {12.8, 9.5, 9.3},
  {14.1, 10.9, 10.2},
  {14.4, 13.8, 12.9},
  {15, 15.1, 16.6},
  {15.2, 15.7, 18.9},
  {15.3, 16.3, 19.3},
  {14.3, 16.7, 17.7},
  {12.1, 14.4, 14.9},
  {10.1, 11.9, 12.4},
  {9.1, 11, 10.7},
  {8.4, 10.2, 9.3},
  {7.6, 9.6, 8.5},
  {8, 9.4, 8},
  {8, 9, 8.2},
  {7.6, 8.8, 8.6},
  {7.5, 8.4, 8.5},
  {7.5, 8.7, 8.2},
  {7, 8.6, 7.8},
  {6.8, 7.9, 7.6},
  {6.9, 7.7, 7.2},
  {6.3, 7.5, 6.9},
  {6.4, 7.3, 6.6},
  {6.6, 7.7, 6.4},
  {9.1, 7.7, 6.4},
  {12.8, 8.7, 6.4},
  {14.4, 10.1, 7.8},
  {15.5, 12.4, 11.6},
  {16, 14.9, 16.3},
  {16.1, 15.8, 18.9},
  {16.7, 17.1, 20.2},
  {15.9, 17, 19.1},
  {12.3, 14.7, 15.4},
  {9.5, 11.6, 12.3},
  {8.4, 10.5, 10.1},
  {7.9, 9.9, 8.8},
  {7.6, 9.5, 7.8},
  {7.4, 9.1, 7.1},
  {7, 9.1, 6.4},
  {7, 8.8, 5.8},
  {6.8, 8.7, 5.4},
  {7, 8.3, 4.9},
  {6.7, 7.9, 4.5},
  {6.1, 7.4, 4},
  {5.9, 7.1, 3.7},
  {5.5, 6.7, 3.6},
  {5.8, 6.6, 3.7},
  {5.9, 6.3, 3.7},
  {7.8, 6.4, 3.6},
  {12.2, 7.1, 5.3},
  {13.8, 10.6, 8.5},
  {14.5, 12.4, 12.8},
  {14.5, 13.5, 16.6},
  {14.7, 14.6, 18.5},
  {14.6, 15.4, 18.5},
  {13.8, 15.2, 16.5},
  {12, 12.9, 13.8},
  {10.4, 11, 11.3},
  {9.6, 10.2, 9.4},
  {8.5, 9.4, 8.3},
  {7.2, 8.6, 7.4},
  {6.7, 8.1, 7.8},
  {5.9, 7.7, 8},
  {5.9, 7.2, 7.8},
  {5.4, 7, 7.3},
  {5.3, 6.5, 7.1},
  {5.6, 6, 6.9},
  {5.5, 6, 6.5},
  {5.6, 5.9, 6.2},
  {5, 5.8, 6.1},
  {4.9, 5.6, 5.7},
  {4.8, 5.3, 5.6},
  {6.6, 5.2, 5.5},
  {9.1, 5.7, 5.9},
  {9.1, 8.2, 6.7},
  {9.6, 9.5, 7.8},
  {9.6, 11, 11.6},
  {9.8, 11.8, 13.4},
  {9, 12.4, 12.5},
  {8.1, 11.2, 11.7},
  {7.3, 9.5, 10.9},
  {7.3, 9, 10.7},
  {7.4, 9.2, 10.8},
  {7.5, 9.4, 10.7},
  {7.4, 9.3, 10.2},
  {7.4, 9.2, 10},
  {7.4, 9, 9.9},
  {7.4, 8.9, 9.8},
  {7.3, 8.7, 9.7},
  {7.3, 8.7, 9.7},
  {7.3, 8.6, 9.7},
  {7.2, 8.7, 9.5},
  {7, 8.6, 9.5},
  {6.9, 8.2, 9.5},
  {7, 8.1, 9.4},
  {7, 8.2, 9.4},
  {7.4, 8.5, 9.7},
  {7.6, 9.2, 10.1},
  {7.7, 9.3, 10.9},
  {7.5, 9.4, 11.4},
  {7.8, 9.5, 11.1},
  {8.1, 9.1, 10.2},
  {8.7, 8.6, 9.9},
  {9.5, 8.6, 10.3},
  {9.1, 8.6, 10.2},
  {8.3, 8.2, 9.9},
  {8.2, 8.4, 9.9},
  {8.2, 8.5, 9.9},
  {8.2, 8.5, 9.9},
  {8.2, 8.6, 9.8},
  {8.2, 8.4, 9.8},
  {7.9, 8.2, 9.8},
  {8, 7.5, 9.6},
  {7.8, 7.1, 9.6},
  {6.2, 6.8, 9.5},
  {5.8, 7, 9.5},
  {5.8, 6.5, 9.6},
  {5.2, 6.5, 9.4},
  {5.3, 6.5, 9.2},
  {6.1, 6.7, 8.8},
  {7.7, 7.6, 8.9},
  {8.9, 8.4, 9.6},
  {9.4, 8.9, 10.6},
  {9.9, 10.2, 11.5},
  {10.2, 10.8, 12.5},
  {11, 11.8, 13.7},
  {11.4, 12.9, 15.8},
  {11.7, 13.5, 16},
  {9, 11.3, 12.9},
  {8, 9.8, 10.9},
  {7.7, 9, 9.6},
  {7.3, 8.7, 8.7},
  {7.4, 8.5, 8.1},
  {7.4, 8.4, 7.6},
  {7.3, 8.1, 7.2},
  {7.1, 8, 6.7},
  {7, 7.7, 6.1},
  {6.7, 7.6, 5.9},
  {6.5, 7.7, 6.4},
  {6.7, 7.8, 7},
  {7.4, 7.8, 7},
  {7.2, 7.9, 6.8},
  {6.2, 7.6, 6.6},
  {6.5, 7.2, 6.5},
  {8.1, 7.7, 6.3},
  {10.8, 8.6, 7},
  {10.9, 10.6, 8},
  {11.1, 9.8, 8.9},
  {11.1, 9.1, 10.3},
  {13, 10.1, 12.9},
  {13, 12.4, 16.1},
  {12.8, 13.7, 16.1},
  {9.4, 11.5, 12.7},
  {7.8, 10.2, 11.6},
  {7.2, 9.3, 9.4},
  {6.8, 8.5, 8.3},
  {6.8, 8.1, 7.3},
  {6.6, 7.8, 6.6},
  {6.9, 7.8, 6.1},
  {6.5, 7.6, 5.6},
  {6.7, 7.4, 5.4},
  {7, 7, 5.2},
  {6.7, 7, 5},
  {6.2, 6.8, 5},
  {5.5, 6.5, 5.1},
  {5.6, 6.3, 5.3},
  {5.3, 6, 5.1},
  {5.5, 6, 5.2},
  {6.7, 6.4, 5.1},
  {10.1, 7, 5.7},
  {10.9, 9, 7.2},
  {11.5, 10.9, 9.8},
  {12, 12.1, 13.8},
  {11.6, 12.3, 14.9},
  {10.2, 11.9, 13.6},
  {9.8, 11.5, 13.2},
  {9.4, 10.5, 12.2},
  {8.7, 10, 11.4},
  {8.5, 9.6, 11.2},
  {8.1, 9.2, 11},
  {7.1, 9.4, 11},
  {7.8, 9.1, 11},
  {8.1, 9.4, 10.8},
  {8, 9.3, 10.5},
  {8.1, 9.2, 10.3},
  {8, 9.2, 10.3},
  {7.9, 9.2, 10.3},
  {7.9, 9.1, 10.2},
  {7.9, 9.1, 10.1},
  {7.9, 9.3, 10},
  {7.9, 9.2, 10},
  {7.9, 9.1, 9.7},
  {7.9, 9.1, 9.8},
  {8, 9.4, 10.1},
  {8.6, 9.5, 10.3},
  {9.1, 10.1, 10.6},
  {9.2, 10.8, 11},
  {8.8, 10.8, 11.3},
  {8.9, 10.6, 11.6},
  {8.7, 10.2, 11.5},
  {8.5, 9.4, 11.3},
  {8.6, 9.2, 10.9},
  {8.5, 9.1, 10.7},
  {8.4, 9.2, 10.7},
  {8.4, 9.3, 10.6},
  {8.1, 9.5, 10.5},
  {7.8, 9.2, 10.4},
  {7.6, 8.7, 10.4},
  {7.5, 8.5, 10.3},
  {7.5, 8.3, 10.2},
  {7.2, 8, 10},
  {7, 7.8, 9.8},
  {6.9, 7.7, 9.4},
  {6.7, 7.5, 9},
  {6.6, 7.5, 9},
  {6.7, 7.4, 9},
  {7.2, 7.4, 8.9},
  {7.4, 7.4, 9},
  {7.2, 7.4, 9.2},
  {7.4, 7.5, 9.4},
  {7.3, 7.5, 9.5},
  {7, 7.6, 9.4},
  {7, 7.7, 9.4},
  {7.2, 7.7, 9.5},
  {7, 7.6, 9.5},
  {7.1, 7.6, 9.4},
  {7.1, 7.6, 9.3},
  {7.4, 7.7, 9.2},
  {7.5, 7.7, 9.1},
  {7.4, 7.7, 9.1},
  {7.2, 7.7, 9.1},
  {7.3, 7.8, 9},
  {7, 7.9, 8.9},
  {6.8, 8, 8.9},
  {6.7, 7.8, 8.8},
  {6.6, 7.6, 8.9},
  {6.6, 7.6, 8.8},
  {6.3, 7.5, 8.7},
  {6.6, 7.5, 8.7},
  {6.8, 7.5, 8.5},
  {7, 7.9, 8.3},
  {8.5, 8.2, 8.5},
  {9.4, 9.5, 9},
  {10.4, 10.6, 9.8},
  {11.2, 12.1, 11.7},
  {12, 12.3, 14.4},
  {12.3, 13.3, 16.7},
  {12.2, 13.4, 15.2},
  {9.4, 11, 12.6},
  {7.7, 9.2, 10.7},
  {7.1, 8.9, 9.3},
  {6.9, 8.4, 8.5},
  {7, 8.4, 7.6},
  {6.5, 8.3, 7.1},
  {6.2, 7.7, 7.2},
  {5.8, 7.5, 7.4},
  {5.7, 7.3, 7.7},
  {6.3, 6.9, 7.6},
  {6, 6.5, 7.5},
  {5.9, 6.5, 7.3},
  {4.9, 6.5, 6.9},
  {4.6, 6.7, 6.6},
  {4.2, 6.2, 6.2},
  {4.8, 5.8, 5.8},
  {6.2, 6.2, 5.7},
  {9, 6.9, 6},
  {9.5, 8.9, 6.3},
  {11.5, 10, 7.9},
  {12.5, 10.4, 10.4},
  {13.1, 11.7, 14.6},
  {12.7, 12.3, 16.5},
  {12.4, 12.9, 15.3},
  {9.9, 10.3, 11.7},
  {8.3, 8.8, 9.6},
  {7.2, 8, 8.2},
  {6.8, 7.5, 7.3},
  {6.4, 7.2, 6.6},
  {6.1, 7, 6},
  {5.9, 7, 5.4},
  {5.8, 7, 4.9},
  {5.6, 6.6, 4.4},
  {5.3, 6.2, 4},
  {5.1, 5.8, 4.2},
  {5.2, 5.4, 4.4},
  {5, 5.2, 4.4},
  {4.6, 4.8, 4.4},
  {4.1, 4.8, 4.3},
  {4.1, 4.5, 4.1},
  {5.4, 4.8, 4},
  {8.6, 5.8, 4.1},
  {10.2, 7.9, 5.1},
  {10.8, 9.3, 7.3},
  {12, 10.5, 11.5},
  {12.1, 11.4, 14.9},
  {11.8, 12.1, 16.1},
  {11.8, 12.6, 14.3},
  {8.5, 9.9, 11.3},
  {6.4, 8.1, 9},
  {5.6, 6.9, 7.4},
  {4.8, 6.6, 6.2},
  {4.8, 6.3, 5.5},
  {4.7, 6.5, 4.7},
  {4.4, 6.2, 4.2},
  {4.5, 6.1, 3.6},
  {5, 6, 3.2},
  {4.2, 5.4, 2.8},
  {4, 5.1, 2.5},
  {3.8, 5, 2.1},
  {3.4, 4.9, 2.6},
  {3.1, 4.9, 2.7},
  {3.5, 4.2, 2.7},
  {3.5, 4.4, 2.7},
  {5.1, 4.9, 2.6},
  {9, 5.8, 3},
  {11, 8.4, 4.8},
  {11.8, 11, 8},
  {12.9, 10.8, 11.9},
  {13.4, 11.2, 13.5},
  {12.7, 12.5, 14.9},
  {12, 12.9, 14},
  {8.5, 10.1, 9.8},
  {8.6, 8.3, 7.9},
  {8.1, 7.7, 6.5},
  {8.1, 7.3, 5.4},
  {6.7, 7.4, 4.5},
  {6.7, 7.6, 3.9},
  {6, 6.8, 3.4},
  {7.1, 6.9, 2.8},
  {5.5, 6.6, 2.4},
  {5.6, 6.2, 1.9},
  {5.2, 6, 1.6},
  {5.3, 5.7, 1.2},
  {3.8, 5.4, 0.9},
  {3.7, 5.3, 0.7},
  {4.4, 5.1, 0.5},
  {4.2, 4.9, 0.4},
  {5.2, 4.9, 0.7},
  {8.9, 6, 1.9},
  {10.8, 7.8, 5.3},
  {12.9, 9.4, 9.4},
  {13.2, 10.9, 13.3},
  {13.4, 11.8, 15.2},
  {12.6, 12.4, 16.6},
  {12.4, 12.8, 14.8},
  {9.1, 10.2, 10.8},
  {6.1, 8, 8},
  {5.7, 7.1, 6.3},
  {5.2, 6.4, 5},
  {4.7, 6, 4.1},
  {4.4, 5.9, 3.3},
  {4.1, 5.5, 2.7},
  {3.6, 5.1, 2.3},
  {3.1, 5, 1.7},
  {3.3, 5.1, 1.3},
  {3.2, 4.9, 0.9},
  {2.8, 4.6, 0.6},
  {2.5, 4.3, 0.4},
  {2.7, 3.9, 0.2},
  {2, 3.9, 0},
  {2.2, 3.4, 0},
  {3.2, 3.6, 0},
  {7.6, 3.6, 1.1},
  {9.4, 5.5, 4.6},
  {10.1, 8.3, 8.6},
  {10.7, 9.2, 11.8},
  {10.5, 10.1, 13.6},
  {10.1, 10.6, 14.6},
  {9.2, 10.8, 12.3},
  {5.9, 8.2, 9.8},
  {4.9, 6.7, 6.8},
  {4.4, 6, 5.4},
  {4.2, 5, 4.2},
  {3.6, 4.9, 3.3},
  {2.8, 5, 2.6},
  {3.2, 5.2, 2.3},
  {2.6, 4.6, 1.7},
  {2.6, 4.3, 1.5},
  {2.3, 4.4, 1},
  {2.9, 4.3, 0.8},
  {2.6, 3.8, 0.7},
  {2.5, 3.7, 0.3},
  {2.4, 3.5, 0.2},
  {2.1, 3.2, 0.2},
  {2.6, 3.2, 0.1},
  {3.9, 3.9, 0.2},
  {6.6, 5.7, 1.6},
  {8.3, 6.5, 4.1},
  {8.8, 7.1, 8},
  {9.5, 8.8, 10.9},
  {9.7, 10.1, 13},
  {9.2, 10.5, 13.8},
  {7.9, 9.7, 11.6},
  {5.6, 7.5, 9.2},
  {3.7, 6.3, 6.8},
  {3.3, 5.3, 5.4},
  {3.5, 4.9, 4.2},
  {3.4, 4.5, 3.4},
  {3.6, 4.2, 3.2},
  {2.4, 3.9, 3.7},
  {2.6, 3.7, 4.1},
  {2.4, 4, 3.5},
  {2.4, 4, 2.8},
  {2, 3.6, 2.3},
  {1.9, 3.2, 1.8},
  {1.8, 3, 1.3},
  {1.8, 2.8, 0.6},
  {1.4, 2.6, 0.1},
  {1.2, 2.5, -0.1},
  {2.5, 2.5, 0.2},
  {5.3, 3.2, 1},
  {7.1, 5.2, 2.3},
  {7.8, 7.8, 4.9},
  {8.4, 8.4, 8.3},
  {8.6, 9.1, 11.8},
  {8.4, 9.4, 12.3},
  {7.5, 9, 10},
  {4.4, 6.9, 8.3},
  {3.2, 5.4, 6.9},
  {2.8, 4.8, 5},
  {2.6, 4.6, 3.8},
  {2.6, 3.9, 3},
  {3.4, 3.7, 2.4},
  {3.2, 3.5, 2.1},
  {2.7, 3, 2.2},
  {3.5, 3.4, 2.9},
  {3.6, 2.8, 3.2},
  {3.6, 3.5, 3.4},
  {3.6, 3.3, 3.6},
  {3.5, 3.2, 3.9},
  {3.5, 2.9, 3.8},
  {3.2, 2.6, 3.6},
  {3.3, 2.6, 3},
  {3.3, 2.6, 3.2},
  {5, 3.2, 3.9},
  {6, 4.5, 5.8},
  {6, 6.5, 8.2},
  {7.3, 7.1, 9.7},
  {7.2, 8.7, 11.5},
  {7.1, 8.5, 11.5},
  {6.3, 8.6, 10.7},
  {5.1, 6.6, 8.6},
  {3.5, 5.1, 6.5},
  {2.8, 4.6, 5.3},
  {4.2, 4.8, 4.2},
  {4.6, 5.2, 4.1},
  {4.4, 4, 4},
  {4.4, 3.6, 3.4},
  {4.4, 3.8, 3},
  {4.4, 3.6, 3.3},
  {4.4, 3.3, 3.6},
  {3.9, 3.1, 3.1},
  {3, 3.1, 2.6},
  {2.4, 3.4, 2.1},
  {1.8, 3, 1.7},
  {2.2, 2.9, 2},
  {2, 2.9, 1.4},
  {2.9, 3, 1.2},
  {5.6, 3.5, 1.9},
  {5.8, 5.3, 4},
  {6.7, 7.2, 6.9},
  {7, 7.6, 10.2},
  {7.7, 8.1, 11.3},
  {7.1, 8.7, 10.3},
  {5.7, 7.8, 9.3},
  {5.1, 6.7, 8},
  {4.9, 6.7, 7.5},
  {5, 6.3, 7.4},
  {5, 6.3, 7.2},
  {4.8, 6.1, 7.2},
  {4.8, 5.9, 7.2},
  {4.6, 5.8, 7.2},
  {4.3, 5.9, 7},
  {3.8, 5.4, 6.8},
  {2.9, 5.2, 5.7},
  {2.3, 6, 4.6},
  {3.3, 5.8, 3.6},
  {3.8, 5.5, 2.4},
  {3.4, 5.5, 1.8},
  {3.1, 5.1, 1.3},
  {3, 4.9, 0.8},
  {3.2, 5.3, 0.6},
  {5.7, 5.5, 0.9},
  {7, 6.3, 4.5},
  {7.9, 7.4, 10.1},
  {7.8, 8.2, 11.5},
  {7.8, 8.7, 11.6},
  {7.5, 8.8, 11.7},
  {7.1, 8.2, 10.7},
  {3.3, 5.9, 6.8},
  {2.3, 4.9, 4},
  {1.3, 4.3, 2.4},
  {1.6, 3.9, 1.2},
  {1.5, 3.5, 0.3},
  {0.9, 2.9, -0.2},
  {-0.3, 2.2, -0.8},
  {-1, 1.8, -1.3},
  {-0.5, 1.4, -1.6},
  {-1.3, 1, -2.1},
  {-1.8, 0.5, -2.5},
  {-2.2, 0.2, -2.8},
  {-2.7, 0, -3},
  {-3, -0.4, -3.4},
  {-3, -0.6, -3.6},
  {-3.1, -0.8, -3.7},
  {-1.9, -0.4, -3.7},
  {1.7, 0.5, -2.9},
  {2.8, 2, 0.1},
  {3.7, 4.2, 3.4},
  {4.3, 5.1, 6.6},
  {5.1, 5.9, 9},
  {5.4, 6.1, 8.7},
  {4.5, 4.9, 7.2},
  {2, 3.4, 4.6},
  {-0.5, 2.6, 2.6},
  {-1.4, 2.5, 1},
  {-1.4, 2.2, -0.3},
  {-1.8, 2.2, -1.1},
  {-1.6, 1.5, -1.8},
  {-1.4, 0.6, -2.3},
  {-1.4, 0.2, -2.6},
  {-2, 0.4, -3.2},
  {-1.9, 0.2, -3.4},
  {-1.6, -0.5, -3.8},
  {-1.7, -0.7, -4.1},
  {-2.4, -0.6, -4.5},
  {-3.3, -0.6, -4.8},
  {-3.8, -0.8, -5.1},
  {-3.5, -0.6, -5.2},
  {-2.9, -0.3, -5.1},
  {0.4, 0.3, -4.1},
  {2, 1.8, -0.9},
  {2.7, 3.5, 2.8},
  {3.1, 4.2, 5.8},
  {3.4, 4.8, 7.3},
  {3.3, 5.1, 7.6},
  {2.7, 4.6, 6.3},
  {0.1, 2.3, 2.3},
  {-1.4, 0.9, 0.2},
  {-2.9, 0.2, -1},
  {-3, -0.1, -2.2},
  {-3.6, -0.6, -2.7},
  {-3.1, -0.9, -3.3},
  {-3.3, -0.8, -3.6},
  {-3.8, -0.9, -4.1},
  {-4, -1.5, -4.6},
  {-5, -1.8, -5},
  {-5.4, -2.3, -5.2},
  {-5.5, -2.2, -5.5},
  {-5.6, -2.5, -5.7},
  {-5.6, -2.8, -6.1},
  {-5.7, -2.9, -6.3},
  {-5.7, -3, -6.4},
  {-4.4, -3, -6.3},
  {-0.8, -2.1, -5.3},
  {1.6, -1.4, -1.4},
  {2.5, 1.8, 1.4},
  {3.2, 2.4, 4.4},
  {4, 3.3, 6.3},
  {4.3, 3.5, 7.1},
  {3.7, 4.1, 5.3},
  {-0.4, 1.3, 1.6},
  {-1.6, 0.2, -0.4},
  {-2, -0.2, -1.5},
  {-2.6, -0.5, -2.3},
  {-2.8, -0.6, -2.8},
  {-2.6, -0.6, -3.3},
  {-2.8, -0.5, -3.7},
  {-2.6, -0.7, -4.2},
  {-2.3, -0.5, -4.5},
  {-2.5, -0.4, -4.7},
  {-2.4, -0.5, -4.9},
  {-2.1, -1.4, -5.1},
  {-2.3, -1.6, -5.4},
  {-2, -1.6, -5.4},
  {-1.8, -1.2, -5.5},
  {-1.8, -1.2, -5.7},
  {-1.3, -1.6, -5.4},
  {3.2, 0.3, -4.5},
  {5.5, 1.1, -0.5},
  {7, 2.8, 2},
  {7.3, 6.3, 5.6},
  {6.9, 8.6, 7.8},
  {5.4, 7.5, 7},
  {6.9, 7.7, 6.6},
  {2.9, 4.4, 2.9},
  {1.7, 4.4, 1.5},
  {1.3, 4.4, 0.1},
  {2.1, 4.2, -0.5},
  {0.4, 3.6, -1},
  {2.4, 3.6, -1.8},
  {1.3, 3.1, -2.3},
  {0.8, 3.1, -2.4},
  {0.1, 2.5, -2},
  {0, 2.6, -2.4},
  {-0.7, 2.2, -2.6},
  {-0.4, 2.1, -2.6},
  {-0.3, 1.6, -3.1},
  {-0.6, 1.1, -3.2},
  {-1.6, 0.6, -3.3},
  {-1.4, 0.4, -3.5},
  {-1.9, 0.1, -3.7},
  {0.6, 0.5, -3.1},
  {2, 1.5, 0.2},
  {2.6, 3.1, 3.9},
  {3.2, 3.6, 7},
  {2.9, 3.4, 7.9},
  {2.5, 4.7, 7.1},
  {2, 4.7, 5.1},
  {-0.1, 3, 4},
  {-0.6, 2, 2.2},
  {-0.3, 1.7, 0.1},
  {-0.9, 1.1, -0.6},
  {-2.1, 1, -1},
  {-3.4, 0.4, -1.7},
  {-3.8, 0.4, -2.3},
  {-3.8, 0.1, -2.1},
  {-2.4, -0.1, -2},
  {-1.1, 0, -1.9},
  {-2.7, -0.4, -1.5},
  {-2.8, -0.5, -2},
  {-3.2, -0.5, -2.7},
  {-4.1, -0.9, -3.3},
  {-4, -1.5, -3},
  {-4.4, -1.5, -3},
  {-3.6, -1, -3.4},
  {-1.2, -0.4, -2.7},
  {-0.2, 0.5, 2.9},
  {0.3, 2.4, 5.3},
  {1.1, 3.1, 5.9},
  {1.5, 3.7, 5.5},
  {1.7, 3.8, 5.3},
  {0.6, 2.6, 4},
  {-1.8, 1.8, 2.1},
  {-2.4, 0.8, 0},
  {-2.7, 1, -1},
  {-2.7, 1.1, -1.5},
  {-2.5, 0.6, -1.3},
  {-2.6, 0.1, -1.1},
  {-2.2, -0.4, -1.6},
  {-2.4, -0.5, -1.5},
  {-2.8, -0.6, -1.6},
  {-3.1, -0.9, -1.6},
  {-3.1, -1.2, -1.7},
  {-3.5, -1.2, -1.9},
  {-3.8, -1.3, -2},
  {-4.1, -1.6, -2.1},
  {-3.9, -1.9, -2.4},
  {-4.2, -2.5, -2.9},
  {-4.2, -1.9, -3.1},
  {-2.3, -1.5, -1.3},
  {-2.3, -1.1, 0.5},
  {-1.5, -0.2, 2.8},
  {-0.8, 0.9, 2.8},
  {-1.3, 1.4, 2.4},
  {-2.4, 1.3, 1.9},
  {-3, 0, 1.5},
  {-3.5, -1, 0.6},
  {-3.5, -1.5, -0.2},
  {-3.3, -2.1, -1.4},
  {-3.6, -2.4, -1},
  {-3.7, -2.3, -1.2},
  {-3.9, -2.4, -2.2},
  {-5.7, -3.2, -3.2},
  {-5.5, -3.1, -3.8},
  {-5.6, -3.1, -3.9},
  {-4.6, -3.3, -3.2},
  {-4, -4, -2.9},
  {-4.4, -3.9, -2.5},
  {-4.3, -3.9, -2.3},
  {-4.3, -4, -2.2},
  {-4.3, -4.1, -2.4},
  {-4.6, -4.3, -3.2},
  {-4.2, -4.1, -3.3},
  {-4.8, -3.8, -2.4},
  {-4.2, -3.6, -1.7},
  {-4.2, -3.7, -1.9},
  {-4.2, -3.6, -1.7},
  {-4.5, -3.1, -1.7},
  {-3.5, -3.1, -1.6},
  {-3.4, -3.4, -1.6},
  {-3.3, -3.4, -1.7},
  {-3.1, -3.2, -1.8},
  {-2.9, -3.1, -1.8},
  {-2.9, -3.1, -1.9},
  {-2.9, -3.1, -1.9},
  {-3, -3.1, -1.8},
  {-2.8, -3.1, -1.8},
  {-3.1, -3.1, -1.8},
  {-3.3, -2.9, -1.8},
  {-3.6, -2.9, -2},
  {-3.6, -2.8, -2.9},
  {-3.6, -2.7, -3.5},
  {-4.3, -3.2, -4.4},
  {-4.7, -3.4, -4.1},
  {-4.1, -3.4, -4.1},
  {-3.6, -3.2, -4.3},
  {-3.2, -2.6, -3.3},
  {-2.8, -2.3, -2.5},
  {-3.1, -2.4, -1.7},
  {-3, -2.2, -1.4},
  {-2.6, -2.6, -1.4},
  {-2.5, -2.3, -1.1},
  {-2.2, -2.4, -1},
  {-2.1, -2.4, -0.5},
  {-2, -2.4, -0.7},
  {-2.8, -2.3, -0.7},
  {-2.7, -2, -0.8},
  {-2.7, -2.1, -0.7},
  {-2.6, -2.1, -0.8},
  {-2.4, -2, -1.2},
  {-2, -2.2, -2.8},
  {-2.1, -2.2, -2.8},
  {-1.7, -1.8, -1.7},
  {-1.6, -1.7, -1.7},
  {-1.9, -2.2, -1.5},
  {-2, -1.8, -1.5},
  {-2, -1.5, -1.6},
  {-1.8, -1.4, -1.5},
  {-1.7, -1.8, -1.7},
  {-2.8, -2.2, -1.7},
  {-2.9, -1.9, -3.9},
  {-1, -1.2, -3.7},
  {0.1, 0.1, -2.1},
  {0, 0.1, -1.3},
  {-0.3, 1.1, 0.3},
  {1.1, 1.7, 0.8},
  {1.2, 1.3, 1.3},
  {-0.3, 1.3, -0.8},
  {-2, -0.1, -3},
  {-2.4, -0.7, -4.6},
  {-3.4, -1.4, -4.7},
  {-3.5, -1.3, -4.4},
  {-3.4, -1.2, -3.7},
  {-4.5, -1.4, -2.8},
  {-4.4, -1.3, -4.3},
  {-4.9, -1.7, -6.1},
  {-4.6, -1.3, -5.6},
  {-4.4, -1, -5.6},
  {-4.7, -1.3, -4.6},
  {-5.3, -2.2, -5.7},
  {-5.5, -2.8, -4.9},
  {-5.8, -3.2, -4.1},
  {-5.9, -3.8, -4.6},
  {-5.8, -4.1, -5.4},
  {-5.6, -4.2, -5},
  {-2.9, -3.9, -4.7},
  {-1, -2.6, -4.3},
  {1, -0.8, -3.3},
  {0.8, 1.2, -1.6},
  {1.9, 1.8, -1},
  {1.1, 1.5, -0.2},
  {-0.5, 0, -1.6},
  {-2.5, -1.4, -3.8},
  {-3.6, -2.2, -5.4},
  {-4.1, -2.8, -6.1},
  {-3.6, -3, -7},
  {-3.6, -3.2, -6.4},
  {-3.5, -3.6, -7.8},
  {-4, -3.6, -8.4},
  {-3.6, -3.9, -9.1},
  {-3.3, -4.2, -9.3},
  {-2.5, -4.1, -7.9},
  {-2.3, -4.2, -6.8},
  {-2.2, -4.4, -7},
  {-2.1, -4.3, -6.1},
  {-2.4, -3.7, -5},
  {-2.9, -3.7, -4.3},
  {-3, -4.3, -4},
  {-2.4, -4.7, -3.6},
  {-1.8, -3.6, -3.2},
  {-1.1, -3.1, -2.5},
  {-2.2, -3.8, -2},
  {-2.1, -3.8, -1.8},
  {-2.4, -3.4, -1.6},
  {-1.6, -3.2, -1.4},
  {-1.2, -2.7, -1.2},
  {-1, -2.8, -1.2},
  {-1.2, -2.6, -1.2},
  {-1.3, -2.3, -1.4},
  {-2, -2.1, -1.8},
  {-2.6, -2.1, -2.9},
  {-2.6, -1.9, -4.2},
  {-3, -1.7, -4.2},
  {-2.6, -1.8, -4.6},
  {-3.1, -2.1, -3.6},
  {-3.5, -2.2, -3.1},
  {-4, -2.3, -3.1},
  {-4, -3.2, -3.4},
  {-4.4, -3.5, -3.3},
  {-4.7, -3.7, -3.3},
  {-4.6, -3.2, -3.8},
  {-4.6, -3.7, -4.4},
  {-4.6, -3.8, -4.7},
  {-2, -3, -4.4},
  {-0.5, -1.7, -3.1},
  {0, 0.5, -2.3},
  {0.4, 0.8, -0.8},
  {1.4, 1.9, -0.3},
  {0.6, 2.4, -1},
  {0.6, 1.8, -2.9},
  {0.1, -0.2, -4.9},
  {0.9, -0.4, -6.2},
  {1, -0.4, -6.6},
  {0.9, -0.5, -7.1},
  {-0.4, -0.6, -6},
  {-0.4, -1, -5.8},
  {-0.7, -1.1, -5.6},
  {-1.2, -1.2, -5.1},
  {-1.6, -1.5, -5},
  {-1.8, -1.6, -4.8},
  {-2.7, -1.8, -4.8},
  {-4.1, -2.3, -5.4},
  {-4.3, -2.6, -5.8},
  {-4.4, -2.6, -6.8},
  {-4.9, -3.2, -7.7},
  {-4.4, -3.3, -7.5},
  {-4.7, -3.4, -9.7},
  {-2.4, -3, -10.5},
  {0, -2.1, -7},
  {1.4, -0.3, -4.7},
  {1.4, 0.7, -2.4},
  {2.6, 1.5, -1},
  {2.2, 1.7, -0.6},
  {1, 1.5, -2.2},
  {-2.4, -1.1, -5.4},
  {-2.9, -1.7, -6.7},
  {-3.7, -2.3, -7.5},
  {-3.8, -2.6, -8.6},
  {-3.2, -3, -8.9},
  {-4.3, -3.2, -9.9},
  {-4.8, -3.3, -10.3},
  {-5.1, -3.5, -10.5},
  {-5.3, -3.9, -10.5},
  {-5.1, -4.1, -10.7},
  {-5.6, -4.4, -11.7},
  {-5.5, -4.4, -11.3},
  {-5.4, -4.5, -11.6},
  {-5.8, -4.8, -9.8},
  {-5.7, -4.9, -9.5},
  {-5.9, -5, -10.6},
  {-5.9, -4.7, -10.9},
  {-3.3, -4.3, -11.7},
  {-3, -3.6, -8},
  {-1.2, -2, -6.7},
  {0.1, -2.4, -4.6},
  {0.7, -2.1, -3.4},
  {0, -1.4, -2.8},
  {-0.7, -1.5, -2.5},
  {0, -2, -2.4},
  {0.4, -2.4, -2.2},
  {0.4, -2.3, -2.1},
  {0.3, -2.1, -2},
  {1, -2, -1.9},
  {1.8, -2, -1.8},
  {1.8, -1.8, -1.7},
  {2.1, -1.7, -1.4},
  {2.2, -1.5, -1.1},
  {1.9, -1.4, -0.5},
  {1.2, -1.1, 0},
  {1.2, -0.9, 0},
  {0.2, -0.9, -0.3},
  {0.2, -0.4, -0.3},
  {0.1, -0.5, -0.3},
  {0.2, -0.4, -0.2},
  {1.5, -0.2, -0.2},
  {2.2, 0, -0.1},
  {1.2, 0.1, 0},
  {1, 0.2, 0.1},
  {2, 0.5, 0.7},
  {2.8, 0.6, 0.8},
  {3.7, 0.3, 0.8},
  {4.2, 0.5, 0.3},
  {2.3, 0.6, 0},
  {1.2, 0.7, -0.1},
  {0.9, 0.4, 0},
  {0.6, 0.5, -0.1},
  {0.5, 0.7, -0.3},
  {0.4, 0.5, 0.1},
  {-0.1, 0.6, 0},
  {0, 0.4, -0.1},
  {-0.1, 0.5, -0.1},
  {-0.3, 0.1, -0.1},
  {-0.1, 0.6, -0.1},
  {0.3, 0.2, -0.3},
  {0.2, -0.1, -0.4},
  {0.1, -0.1, -0.4},
  {-0.2, -0.4, -0.4},
  {-1, -0.1, -0.5},
  {-1.2, -1, -0.7},
  {0.5, -0.6, -0.9},
  {2.9, -0.3, -1.2},
  {4.3, 0.2, -1.2},
  {5.1, 1.8, -0.8},
  {4.9, 1.2, -0.5},
  {4.2, 1.4, -0.1},
  {3.3, 1.1, 0},
  {2.5, 0.6, -0.1},
  {2.2, 0.8, 0},
  {2.3, 0.6, 0},
  {2.3, 0.2, 0},
  {2.5, 0.3, 0},
  {2.6, 0.2, 0},
  {2.4, 0.2, 0},
  {2.1, 0.5, 0},
  {1.5, 0.4, 0},
  {1.2, 0.1, 0.2},
  {1.3, 0.3, 0.1},
  {1.6, 0.1, 0.1},
  {1.3, 0.3, 0.1},
  {0.6, 0, 0},
  {0.7, 0, -0.2},
  {1, 0, -0.2},
  {1.3, 0.1, -0.2},
  {1.6, 0.3, 0.2},
  {1.8, 0.6, 0.9},
  {3.1, 1.1, 1.3},
  {4.2, 1.9, 2.2},
  {3.9, 2.4, 3.1},
  {2.6, 2.1, 2.3},
  {2.1, 1.6, 2},
  {1.9, 1.2, 1.2},
  {2.4, 0.9, 0.7},
  {2, 0.7, 0.1},
  {2.1, 0.7, 0.2},
  {1.6, 0.7, 0.5},
  {1.5, 0.8, 0.4},
  {1.4, 0.7, 0.4},
  {0.6, 0.5, 0.3},
  {-0.2, 0.2, 0.5},
  {-0.3, 0.5, 0.5},
  {0.2, -0.1, 0.3},
  {-0.9, 0.3, 0.1},
  {-1, 0.6, -0.1},
  {-0.7, 0.8, -0.1},
  {-0.2, 1.1, -0.3},
  {-0.8, 1.1, -0.2},
  {-0.3, 1.2, -0.3},
  {0.8, 1.7, -0.4},
  {1.7, 2.1, -0.1},
  {1.8, 2.1, 0.2},
  {2.7, 1.7, 0.5},
  {2.1, 1.5, 0.7},
  {2, 1.5, 0.8},
  {2.4, 1.6, 1},
  {2.4, 1.2, 0.9},
  {1.7, 1.2, 0.3},
  {1, 1.2, 0},
  {0.7, 1, -0.3},
  {0.7, 0.8, -0.9},
  {-0.1, 0.5, -1.3},
  {-0.2, 0.2, -0.8},
  {-0.9, 0, -0.2},
  {-0.9, 0.6, 0},
  {-1.2, 0.7, -0.1},
  {-1.1, 0.4, -0.4},
  {-0.6, -0.2, -0.8},
  {-0.9, -0.5, -1},
  {-1.5, -0.8, -1.2},
  {-1.3, -0.9, -1.4},
  {-1.6, -1.2, -1.7},
  {-2.1, -1, -2},
  {0.5, -0.4, -2.2},
  {2.8, 0.4, -2.5},
  {2.9, 2, -2.4},
  {3.5, 3.7, -1.1},
  {4.2, 4.1, 1.3},
  {4.1, 4.3, 2.3},
  {3.7, 3.4, 0.8},
  {-0.1, 1.6, -1.7},
  {-0.8, 0.4, -3.9},
  {-1.5, 0, -4.9},
  {-1.7, -0.1, -5.6},
  {-1.9, -0.4, -5.9},
  {-2.4, -0.6, -6.3},
  {-2.8, -1.3, -6.7},
  {-2.8, -1.5, -8},
  {-3.1, -1.7, -8.2},
  {-2.7, -1.6, -8.2},
  {-3.1, -2, -8.5},
  {-4, -2.5, -9.1},
  {-4.1, -3.1, -9.1},
  {-3.8, -3, -9.1},
  {-3.7, -3.2, -8.8},
  {-3.8, -3.4, -9.2},
  {-3.9, -3.2, -9.2},
  {-1.7, -3.2, -9.6},
  {0.4, -2.6, -6.9},
  {1.7, 0.2, -4.8},
  {0.8, -0.6, -3.8},
  {0.7, -0.7, -2.5},
  {0.2, -0.7, -2.1},
  {-0.3, -0.9, -1.9},
  {-1.4, -1, -1.8},
  {-1.5, -1.4, -1.9},
  {-1.4, -1.8, -2},
  {-1, -2, -2.7},
  {-1.5, -1.8, -2.7},
  {-1.8, -1.5, -2.8},
  {-2, -1.5, -2.6},
  {-1.1, -1.6, -2.9},
  {-1.1, -1.6, -3.1},
  {-1.4, -1.6, -3.1},
  {-0.4, -1.9, -3.5},
  {-0.1, -1.7, -3.6},
  {0, -1.7, -4},
  {-0.7, -1.7, -4.3},
  {-0.2, -1.4, -5.2},
  {0.1, -1.1, -5.6},
  {0.4, -1.4, -6.2},
  {1, -1.2, -5.6},
  {1.7, -0.4, -4.1},
  {2.5, 1.2, -1.3},
  {2.8, 2, -0.3},
  {3.6, 2.6, -0.2},
  {3.5, 4, 1.2},
  {3, 4, 0.3},
  {2.2, 2.9, -1.2},
  {1.8, 2.2, -3.1},
  {1.3, 1.6, -4.6},
  {0, 1.2, -5.2},
  {0, 1.2, -6},
  {-1.2, 0.5, -6.7},
  {-2.1, 0.3, -7.2},
  {-2.3, 0, -7.1},
  {-2.6, -0.4, -8},
  {-3.4, -0.8, -8.2},
  {-4.2, -1.2, -8.8},
  {-4.1, -1.7, -8.6},
  {-4.5, -1.9, -9.3},
  {-4.6, -2.6, -9.8},
  {-4.9, -3, -10.3},
  {-4.8, -3.2, -10},
  {-5.2, -3.1, -9.6},
  {-2.7, -3.8, -9.1},
  {-0.2, -2.5, -6.7},
  {0, -0.5, -5},
  {0.9, 0.9, -2.2},
  {1.5, 1.4, 0.2},
  {1.2, 1.7, 0.8},
  {0.8, 0.7, -0.8},
  {-3.2, -1, -3.9},
  {-4.2, -1.6, -5.9},
  {-4.6, -2.2, -6.8},
  {-4.6, -2.9, -7},
  {-4.7, -2.8, -8.5},
  {-4.7, -3, -8.8},
  {-5.2, -3.1, -9.2},
  {-5.6, -3.2, -9.8},
  {-6.2, -3.8, -10.9},
  {-6.5, -4.1, -10},
  {-6.3, -4.4, -10.8},
  {-6.4, -5.1, -11},
  {-6.6, -5.4, -10.9},
  {-6.2, -5.7, -11.7},
  {-6, -5.9, -11.7},
  {-5.8, -5, -11.9},
  {-4.7, -5.6, -12.3},
  {-2.9, -5.1, -11.7},
  {-2.1, -3.6, -9.6},
  {-0.6, -1.5, -6.2},
  {0.7, -0.8, -2.9},
  {1.4, 0.5, -1.4},
  {2.8, 1.2, -0.1},
  {1.6, 0.8, -2},
  {0.4, -0.7, -3.9},
  {-0.5, -0.7, -5.1},
  {-2.2, -0.6, -5.8},
  {0, -2, -7.3},
  {1.3, -1.4, -7.7},
  {1.7, -1.4, -8.2},
  {1.8, -1.1, -8.4},
  {1.8, -0.4, -8.7},
  {1.3, -0.5, -8.3},
  {1.9, -0.7, -7.8},
  {1.4, -0.1, -7.8},
  {1.7, -1.2, -7.9},
  {1.2, -1.3, -7.7},
  {1.2, -1, -7.1},
  {-0.3, -1.4, -6.7},
  {-0.9, -1.2, -6.8},
  {-0.8, -0.9, -6.9},
  {1, -0.5, -6.4},
  {1.6, 0.6, -4.7},
  {1, 2.5, -2.6},
  {2.3, 1, -1.8},
  {3.3, 1.9, -0.3},
  {3.3, 2.1, 0.1},
  {2.1, 1.3, 0.1},
  {1.5, 1.4, 0.1},
  {2.4, 1.4, 0.1},
  {1.4, 1.3, 0.1},
  {1.2, 1.3, 0.2},
  {0.2, 1.1, 0.2},
  {0.2, 0.5, 0.1},
  {0.8, 0.1, 0},
  {1.8, -0.4, -0.1},
  {1.6, 0.4, -0.1},
  {1.6, 0.5, -0.1},
  {1.4, 0.7, -0.1},
  {1.2, 0.7, -0.1},
  {0.9, 1.5, -0.1},
  {1.1, 1, -0.1},
  {1.3, 1.4, -0.1},
  {1.3, 1.7, -0.1},
  {1.6, 1.5, 0},
  {2.4, 2, 0.3},
  {2.9, 3.3, 1.4},
  {3.5, 4, 2.1},
  {4.5, 4.4, 3},
  {6.7, 5.6, 4.5},
  {6.6, 5.8, 4.6},
  {5, 5.2, 3.3},
  {3.2, 3.5, 1.3},
  {2.2, 2.6, 0},
  {2.5, 2.7, -0.5},
  {2.2, 2.3, -1.5},
  {1.7, 2.2, -1.5},
  {1.9, 2.3, -0.7},
  {0.8, 1.5, -0.1},
  {0.5, 1, 0},
  {0.7, 0.9, 0},
  {0.6, 1.3, 0},
  {0.5, 0.9, -0.1},
  {0.3, 0.2, -0.2},
  {-0.7, 0.5, -0.3},
  {-1, 0.3, -0.4},
  {-1.1, 0.4, -0.4},
  {-1.4, 0.5, -0.6},
  {-1.1, -0.4, -0.8},
  {0.1, 0.2, -0.8},
  {2.7, 2.3, -1.1},
  {4.5, 3.4, -1.2},
  {5.8, 4.3, -1.1},
  {6.4, 5.1, -0.5},
  {5.3, 5.3, -0.4},
  {4.5, 4.9, -0.8},
  {0.7, 3, -1.7},
  {-0.6, 2.5, -2.5},
  {-0.8, 2.1, -3.1},
  {-1.3, 2, -3.3},
  {-1.3, 1.8, -2.9},
  {-1.3, 1.6, -2.6},
  {-1.8, 1, -2.6},
  {-2.1, 0.8, -2.9},
  {-1.5, 0.4, -3.1},
  {-2.2, 0.5, -3.2},
  {-3.1, 0, -3.4},
  {-3.1, -0.2, -3.7},
  {-3.2, -0.4, -4},
  {-4.3, -0.5, -4.4},
  {-4.2, -0.8, -4.5},
  {-4.6, -1.5, -4.9},
  {-4.4, -1.4, -5.7},
  {-2.5, -1.5, -6.8},
  {0.1, -1.2, -5.6},
  {1, 0.7, -3.5},
  {2.2, 1.6, -1.9},
  {2, 1.9, -0.5},
  {2.4, 2.5, -0.2},
  {1.8, 1.4, -1.3},
  {-1.1, 0.1, -3},
  {-1.7, -0.7, -4.3},
  {-2, -1, -5.1},
  {-1.8, -1, -5.8},
  {-1.1, -0.5, -6.4},
  {-0.8, -0.4, -6.7},
  {-0.6, -0.5, -7.1},
  {-1.2, -2.3, -7.1},
  {0, -2.2, -7.1},
  {0.4, -2, -7.5},
  {0.2, -0.7, -7.3},
  {-0.1, 0.5, -7.6},
  {-0.1, 0.7, -7.8},
  {0, 0, -8},
  {-0.1, -0.2, -7.9},
  {-0.3, -0.3, -7.7},
  {0, -0.2, -8},
  {1.8, 0.5, -7.6},
  {2, 0.9, -5.8},
  {3.3, 1, -3.8},
  {3.7, 2.2, -2},
  {2.7, 2.8, -1},
  {2.7, 2.1, -0.7},
  {2.2, 1.3, -1.1},
  {1.3, 0.6, -2.5},
  {1.3, 0, -3.5},
  {1.5, -0.7, -3.6},
  {1.5, -1, -3.8},
  {1.4, -0.8, -4.8},
  {1.5, -0.2, -5.1},
  {2.3, 2, -5.4},
  {3.1, 5.4, -5.4},
  {2.6, 4.2, -5.3},
  {2.6, 4, -5.7},
  {1.7, 4.6, -5.8},
  {1.3, 4.8, -4.7},
  {1.3, 3.3, -4.2},
  {0.6, 2.7, -4},
  {0.2, 2.3, -4.4},
  {-0.5, 1.7, -4},
  {0.3, 1.5, -4.7},
  {1, 2.3, -4.7},
  {3.5, 2.8, -3.2},
  {4.2, 4.3, 0},
  {4.3, 4.4, 5.1},
  {3.1, 2.9, 7.3},
  {2.6, 2.1, 6.2},
  {1.2, 0.2, 5.3},
  {-0.4, -0.2, 3.4},
  {-1.5, -0.5, 2.6},
  {-2.3, -1, 1.1},
  {-2.5, -1.1, -0.7},
  {-3.1, -1.7, -1.6},
  {-5.3, -2.1, -2.7},
  {-6, -2.2, -3.9},
  {-5.5, -2.5, -4.4},
  {-5.4, -2.6, -4.1},
  {-5.6, -2.6, -4.7},
  {-4.5, -3.1, -4.6},
  {-4.9, -3.5, -4.6},
  {-6.6, -3.8, -6.4},
  {-6.3, -3.5, -7.1},
  {-4.6, -3.2, -8.4},
  {-4.7, -3.8, -8.8},
  {-4.3, -3.6, -9.4},
  {-2.8, -2.3, -9},
  {-1.5, -1.8, -7.3},
  {-0.6, -0.2, -4.3},
  {-0.2, 0.5, -1.1},
  {-0.2, 1.2, 1.4},
  {-0.3, 1, 1.8},
  {-0.8, 0.5, 0.3},
  {-2.9, -0.7, -3.1},
  {-4.9, -1.2, -4.8},
  {-5.8, -1.9, -6.4},
  {-5.6, -2.8, -8.1},
  {-5.2, -3.2, -8.9},
  {-5.4, -3.7, -10},
  {-5.3, -3.7, -9.9},
  {-5.1, -4, -10.2},
  {-6.7, -4.6, -11.2},
  {-6.8, -5.2, -12.1},
  {-7.2, -5.6, -12},
  {-7.9, -5.2, -12.2},
  {-7.7, -5.4, -12.7},
  {-7.9, -5.5, -12.8},
  {-7.7, -5.4, -12.7},
  {-7.5, -5.7, -12.9},
  {-7.6, -5.7, -13.2},
  {-5.4, -4.8, -12.9},
  {-2.1, -3.7, -9.4},
  {-2.7, -3.5, -7.6},
  {-2.5, -2.9, -6.5},
  {-2.3, -2.6, -4.7},
  {-1.8, -2.5, -4.1},
  {-1.6, -3.2, -3.9},
  {-3, -2.8, -5.3},
  {-2.9, -3.1, -6.8},
  {-3.4, -3.1, -6.1},
  {-3.2, -2.8, -6.9},
  {-3.7, -2.9, -7.6},
  {-4.1, -3.4, -7.9},
  {-4.1, -3.7, -8},
  {-4.6, -3.5, -9.5},
  {-5, -4, -9.7},
  {-4.8, -3.8, -9.9},
  {-5.1, -3.5, -10.3},
  {-5.1, -4.2, -10.7},
  {-5.4, -4.5, -11.2},
  {-5.4, -4.9, -11.4},
  {-5.6, -5.2, -11.8},
  {-5.1, -5, -11.9},
  {-4.5, -3, -11.7},
  {-2.1, -3.6, -11.4},
  {1, -3.6, -8.5},
  {3.1, -1.2, -4.8},
  {3.8, 1.9, -1.7},
  {2.9, 2.8, -0.5},
  {2.9, 0.6, -0.1},
  {2.4, 0.9, -0.7},
  {0.2, -0.1, -2.3},
  {-0.9, -0.7, -3.4},
  {-0.7, -0.7, -3.5},
  {-1.4, -1.2, -5.2},
  {-2, -1.5, -6.5},
  {-1.7, -1.4, -7.5},
  {-2.7, -1.6, -8.1},
  {-3.3, -1.9, -8.5},
  {-3.1, -2.2, -8.8},
  {-3.2, -1.7, -9.2},
  {-3.7, -2.2, -9.4},
  {-3.9, -2.4, -9.8},
  {-3.5, -3.3, -10.6},
  {-3.3, -2.6, -10.3},
  {-3.6, -3.5, -10.4},
  {-3.1, -3, -11},
  {-1.9, -3.5, -11.1},
  {-0.2, -2.2, -10.9},
  {3.5, -1.9, -9},
  {4.6, 0.9, -5},
  {5.2, 3.2, -1.9},
  {5.3, 3.7, 0.5},
  {5.4, 3.9, 1.4},
  {4.5, 2.9, -0.6},
  {-0.1, 0.7, -3.5},
  {-1.4, -0.2, -5.3},
  {-1.2, -0.5, -6.4},
  {-1.6, -0.6, -7.1},
  {-1.6, -0.9, -7.9},
  {-2, -0.9, -8.7},
  {-2.3, -1.1, -9.2},
  {-2.5, -1.3, -8.8},
  {-3.4, -1.3, -9.7},
  {-3.1, -1.8, -9.8},
  {-3.6, -1.9, -10.4},
  {-3.5, -2.1, -10.4},
  {-3, -1.9, -10.5},
  {-3, -2.1, -9.8},
  {-3.4, -2.6, -10.6},
  {-4.1, -2.8, -10.5},
  {-3.2, -2.4, -10.9},
  {-2.5, -2.6, -10.6},
  {-0.3, -3, -8.6},
  {2, -1.4, -5.3},
  {2.2, -0.9, -3.2},
  {2.7, 0.6, -1.5},
  {2.9, 0.5, -0.4},
  {2.2, -0.1, -1.7},
  {-0.7, -0.5, -3.8},
  {-1.5, -0.9, -5.4},
  {-1.8, -1.2, -5.7},
  {-2.2, -1.3, -6.7},
  {-2.5, -1.6, -7.4},
  {-2.1, -1.7, -7.8},
  {-1.4, -1.5, -8.3},
  {-1, -1.5, -8.4},
  {-1.2, -1.5, -9},
  {-1.3, -1.5, -9},
  {-1.5, -1.6, -8.8},
  {-1.6, -1.9, -9},
  {-1.8, -2, -9.5},
  {-1.8, -1.9, -9.8},
  {-1.6, -1.9, -10},
  {-1.9, -2.1, -10.1},
  {-1.3, -1.9, -9.6},
  {0.3, -1.3, -9.5},
  {2.2, -0.6, -7},
  {4.1, 1.7, -3.5},
  {4.3, 3.4, -0.1},
  {4.8, 4.8, 2},
  {5, 4.7, 3.1},
  {3.8, 2.7, 0.9},
  {0.6, 1.5, -1.9},
  {-0.4, 1.3, -3.2},
  {-1, 0.1, -4.8},
  {-1.5, -0.1, -5.7},
  {-1.4, -0.4, -6.3},
  {-2.1, -0.8, -6.9},
  {-2.6, -1, -7.2},
  {-2.2, -1.2, -7.6},
  {-2.4, -1.3, -8},
  {-2.5, -1.5, -8.1},
  {-2.7, -1.5, -8.6},
  {-3, -1.6, -8.5},
  {-3.3, -1.8, -9.1},
  {-2.8, -1.8, -8.8},
  {-3.2, -1.5, -8.9},
  {-2.9, -2, -9.8},
  {-2.8, -2, -9.5},
  {-0.8, -1.8, -9.5},
  {1.9, -1.3, -7.2},
  {3.8, 1.6, -3.6},
  {4.8, 3.9, -1.1},
  {5, 4.5, 1.9},
  {4.7, 4, 2.7},
  {4.5, 3.7, 0.7},
  {1.8, 1.6, -1.7},
  {-0.6, 0.5, -3.4},
  {-0.2, 0, -4.4},
  {0.6, -0.2, -5.2},
  {0.3, -0.6, -6},
  {0.1, -0.8, -6.7},
  {0.6, -1.1, -6.7},
  {0.8, -1.2, -7.4},
  {0.6, -1.2, -7.3},
  {-0.2, -1.5, -7},
  {-0.6, -1.7, -7.5},
  {-0.5, -1.8, -8},
  {-1.4, -2.1, -7.7},
  {-2.1, -2.2, -8.3},
  {-2.1, -2, -8},
  {-1.9, -1.9, -7.2},
  {-1.4, -1.1, -7.1},
  {-0.5, -0.9, -6.2},
  {0.3, -0.3, -4.7},
  {1.1, 0.3, -3.5},
  {1.8, -0.2, -1.6},
  {2.4, 0.1, -0.5},
  {2, 0.9, 0.4},
  {0.4, 0.9, -0.2},
  {-0.1, -0.2, -2.4},
  {-0.5, -0.9, -2.7},
  {-0.6, -0.6, -5},
  {-0.9, -0.8, -5.7},
  {-1.6, -0.9, -6.4},
  {-1.7, -1.1, -7.4},
  {-2.2, -1.5, -7.6},
  {-1.9, -1.6, -7.8},
  {-2.5, -1.9, -8.4},
  {-3, -2, -9.1},
  {-3, -2.1, -9.1},
  {-3.2, -2.6, -9.1},
  {-3.5, -3.1, -9.3},
  {-2.1, -2.7, -9.4},
  {-1.8, -2.8, -8.1},
  {-1.8, -2.5, -6.8},
  {-2, -1.9, -6.3},
  {-1.7, -1.8, -5.4},
  {-1.7, -1.4, -4.3},
  {-1.3, -0.8, -3.2},
  {-1, -0.3, -2.5},
  {-0.7, -1.1, -1.8},
  {-0.1, -0.3, -1.2},
  {0, 0, -1.1},
  {-0.8, -0.7, -1.3},
  {-1, -0.7, -1.7},
  {-1.4, -0.6, -1.7},
  {-1.3, -0.9, -1.4},
  {-1.3, -1.4, -1.4},
  {-1.9, -1.4, -1.6},
  {-1.3, -1.9, -1.8},
  {-1.5, -1.8, -2},
  {-1.8, -1.5, -1.9},
  {-2.8, -1.7, -2},
  {-3, -2.1, -2.2},
  {-3.6, -2.1, -2},
  {-3.7, -2.3, -1.9},
  {-4.2, -2.7, -1.9},
  {-4.2, -3, -1.8},
  {-4.5, -3.5, -1.9},
  {-4.6, -3.3, -1.8},
  {-4.3, -2.7, -2},
  {-4.1, -2.1, -1.4},
  {-3.5, -1.9, -0.8},
  {-3.2, -1.8, -0.6},
  {-3.4, -2.3, -0.5},
  {-3.2, -2.7, -0.4},
  {-3.1, -3.1, -0.9},
  {-3, -2.9, -0.8},
  {-3.2, -2.7, -0.8},
  {-3.5, -2.7, -0.7},
  {-3.8, -2.6, -1.6},
  {-4.2, -2.6, -3.6},
  {-5.5, -2.6, -3.3},
  {-5.3, -2.6, -2.4},
  {-6.2, -2.7, -2.2},
  {-6.2, -3.5, -2.4},
  {-6.3, -3.9, -2.7},
  {-5.6, -4, -2.9},
  {-5.7, -3.9, -3.2},
  {-5.1, -3.9, -3.9},
  {-4.8, -3.6, -4.6},
  {-4.7, -3.7, -4.5},
  {-4.5, -3.7, -4.6},
  {-5, -3.6, -4},
  {-5, -3.6, -3.6},
  {-4.9, -3.4, -3.1},
  {-5.2, -3.2, -2.7},
  {-4.8, -3.4, -2.3},
  {-4.7, -3.2, -1.5},
  {-5, -3.1, -1.4},
  {-5.1, -2.6, -1.4},
  {-5.4, -2.8, -1.5},
  {-5.4, -4.1, -1.5},
  {-5.4, -4.3, -1.6},
  {-5.5, -3.9, -2},
  {-5.9, -3.4, -1.9},
  {-6.1, -3.3, -2.3},
  {-6.3, -3.7, -2.5},
  {-6.5, -3.4, -2.8},
  {-6.8, -3.4, -4.2},
  {-7.1, -3.6, -5},
  {-7.4, -3.7, -4.8},
  {-7.4, -3.7, -5.2},
  {-7.5, -3.8, -5.8},
  {-7.3, -3.9, -5.9},
  {-7, -3.9, -6.7},
  {-7.1, -4, -6.9},
  {-7, -4.1, -7.5},
  {-6.1, -4.1, -6.6},
  {-5.4, -4, -5.6},
  {-4.1, -3.7, -4.8},
  {-3.2, -3.4, -3.4},
  {-3.4, -2.8, -2.6},
  {-3.9, -2.1, -3.2},
  {-5.5, -2.6, -5.1},
  {-7.9, -3.8, -7.6},
  {-8.8, -4.6, -9.7},
  {-9.3, -5.2, -10.9},
  {-9.5, -5.5, -12.2},
  {-10, -6, -13.5},
  {-9.9, -6.4, -13.9},
  {-10.2, -6.8, -14.6},
  {-10.7, -7, -15.7},
  {-10.9, -7.5, -16.1},
  {-11, -7.8, -17},
  {-11.7, -8.2, -16.9},
  {-11.4, -8.3, -17.1},
  {-11.3, -8.6, -17.5},
  {-11.6, -8.8, -17.6},
  {-11.9, -9.3, -17.5},
  {-12, -9.3, -18.2},
  {-11.5, -9.4, -18.9},
  {-10.7, -9.4, -18.2},
  {-8.6, -8.1, -14.8},
  {-5.8, -7.1, -10.3},
  {-5.4, -6, -8.2},
  {-4.8, -4.8, -6.6},
  {-5.2, -4.3, -6.5},
  {-6.7, -4.8, -8.3},
  {-8.4, -6.2, -11.2},
  {-9.6, -7.1, -13.5},
  {-9.7, -7.6, -13.6},
  {-9.9, -7.9, -14.4},
  {-9.9, -8.3, -14.7},
  {-9.5, -8.4, -15.1},
  {-7.7, -7.7, -13.3},
  {-7, -7.4, -11.1},
  {-7.5, -6.9, -10.7},
  {-8.6, -7.4, -12},
  {-9.5, -7.9, -13.1},
  {-9.4, -8.2, -13.4},
  {-9.1, -8.5, -13.8},
  {-8.6, -7.8, -13.2},
  {-7.9, -7.7, -12.6},
  {-7.7, -7, -12.3},
  {-7.9, -6.9, -13},
  {-7.4, -6.6, -12.7},
  {-6.3, -5.5, -12.6},
  {-5.7, -4.8, -12.2},
  {-4.9, -5.5, -10.8},
  {-4.5, -4.7, -9},
  {-4.1, -4.3, -8.8},
  {-4.6, -4.6, -7.9},
  {-4.6, -4.6, -6.7},
  {-4.7, -4.2, -6},
  {-5.3, -4.5, -5.7},
  {-5, -4.6, -5.4},
  {-4.7, -4.6, -5.2},
  {-4.6, -4.4, -5},
  {-4.8, -3.8, -4.8},
  {-4.8, -4.4, -4.7},
  {-4.6, -4.8, -4.6},
  {-4.5, -5.7, -4.6},
  {-4.2, -5.3, -4.5},
  {-3.5, -5.2, -4.4},
  {-3.3, -4.6, -4.5},
  {-3, -3.6, -4.3},
  {-3.4, -3.1, -4.2},
  {-3.2, -3, -4.1},
  {-3.6, -2.8, -3.9},
  {-3.1, -2.1, -3.5},
  {-2.4, -2, -2.8},
  {-1.8, -1.6, -2.1},
  {-0.9, -0.9, -1.8},
  {-0.6, -0.6, -1.6},
  {-0.4, -1, -1.2},
  {-0.9, -1.4, -1.1},
  {-1.2, -2.2, -1.1},
  {-1.2, -1.8, -1.1},
  {-1.5, -0.6, -1.2},
  {-0.7, -0.1, -1.7},
  {-0.8, 0.2, -2.5},
  {-0.9, 1.4, -3.1},
  {-0.4, 1.4, -3.4},
  {-0.1, 1.4, -3.1},
  {0.2, 1.3, -2.6},
  {-0.8, 1.7, -2.1},
  {-0.7, 1.7, -2},
  {-0.3, 1.5, -2.2},
  {-0.1, 1.4, -2.2},
  {1.4, 1.5, -2},
  {1.9, 1.9, -2},
  {2.2, 2.1, -2.2},
  {2.2, 2, -2.7},
  {2.1, 2.5, -2.1},
  {2.2, 3.1, -1.1},
  {2.4, 3.5, -0.6},
  {2.4, 3.9, 0},
  {2.8, 4.2, 1},
  {3.3, 4.3, 1},
  {2.3, 4.1, 1},
  {1.8, 3.4, 0.1},
  {2.8, 3.7, -0.3},
  {3, 4.1, 0.7},
  {2.9, 3.9, 0.9},
  {3.1, 3.5, 0.4},
  {1.9, 3, -0.4},
  {1.2, 2.9, -0.9},
  {1.8, 2.8, -1.1},
  {2.3, 2.3, -1.4},
  {1.2, 2.6, -1.5},
  {1.2, 3.1, -1.9},
  {1.9, 2.9, -1.9},
  {1.6, 3, -2},
  {0.8, 2.8, -1.9},
  {0.1, 2.7, -3.6},
  {0, 2.8, -3.7},
  {2.3, 3.2, -3.2},
  {1.6, 3.5, -2.6},
  {2.2, 3.7, -1.2},
  {2, 4, -0.1},
  {3.2, 4.5, 1.1},
  {3.3, 4.7, 2.3},
  {3, 4.8, 2.9},
  {2.3, 4.7, 3},
  {1.4, 4.3, 2.8},
  {0.4, 3.8, 1.8},
  {0.1, 3.4, 0.8},
  {1.1, 3.1, -0.6},
  {1.1, 2.5, -0.7},
  {0, 2, -1.3},
  {0.1, 1.6, -3.5},
  {-1.4, 1.4, -4.6},
  {-1.8, 0.8, -5.3},
  {-1.8, 0.5, -6.3},
  {-2.1, 0.2, -7.8},
  {-2.6, -0.5, -8.3},
  {-2.9, -0.8, -8.9},
  {-3, -1.1, -9.5},
  {-3.8, -1.3, -9.6},
  {-4.2, -1.7, -10.5},
  {-4, -2, -10.5},
  {-2.5, -1.7, -10.8},
  {-1.2, -1.3, -8.1},
  {0.7, -0.1, -5},
  {1.5, 1.2, -2.5},
  {1.5, 1.8, 0.2},
  {1.9, 2.3, 1},
  {0.6, 2.3, -0.5},
  {-1.6, 0.4, -3.8},
  {-2.9, -0.7, -5.7},
  {-3.6, -0.8, -7.2},
  {-3.7, -1.2, -7.9},
  {-2.5, -2, -8.8},
  {-2.1, -2.1, -8.9},
  {-1.7, -1.9, -8.7},
  {-2.3, -2.1, -8.4},
  {-1.9, -1.8, -8.3},
  {-1.9, -1.7, -6.4},
  {-2.6, -1.9, -5.8},
  {-2.7, -2.2, -5.5},
  {-2.4, -2.8, -5.1},
  {-2.9, -2.8, -5.8},
  {-2.9, -2.6, -6.7},
  {-2, -2.3, -5.5},
  {-2.3, -2.4, -4.9},
  {-2.2, -2.1, -4.1},
  {-1.2, -1.3, -2.8},
  {-1.3, -0.8, -1.8},
  {-1.2, -0.2, -0.5},
  {-0.9, 0.1, 0.4},
  {-1, 0.5, 0.7},
  {-0.9, 0.7, 0.5},
  {-1, -0.1, -0.1},
  {-1, -0.5, -0.3},
  {-1.1, -0.1, -0.9},
  {-1, -0.2, -1.1},
  {-1.3, -0.6, -1.4},
  {-1.1, -1.1, -1.3},
  {-1.3, -0.9, -1.5},
  {-1.6, -0.8, -1.7},
  {-1.8, -0.9, -1.9},
  {-1.8, -1.3, -2.7},
  {-2.5, -1.8, -3.6},
  {-3.5, -2.1, -5.5},
  {-4.5, -2.5, -7.3},
  {-4.8, -2.9, -7.9},
  {-4.9, -3.3, -8.8},
  {-4.6, -3.3, -9.2},
  {-4.5, -3.4, -9.5},
  {-3.2, -2.8, -10.1},
  {-1.2, -2, -6.9},
  {0.6, -0.4, -3.7},
  {2.6, 0.9, -0.9},
  {2.6, 1.4, 1.2},
  {2.4, 2.8, 2.2},
  {1.8, 2.6, 0.3},
  {-0.8, 0, -2.9},
  {-1.8, -0.5, -5.2},
  {-2.8, -0.6, -5.6},
  {-2.9, -1, -7.4},
  {-2.6, -0.8, -7.3},
  {-1.5, -0.7, -6.2},
  {-1.2, -0.7, -4.5},
  {-0.7, -0.8, -4.4},
  {-0.6, -0.4, -5.1},
  {-0.4, -0.6, -6.1},
  {-0.5, -0.8, -6},
  {-0.4, -1, -5.4},
  {-1.1, -1.2, -5.2},
  {-1.9, -1, -6.8},
  {-2.3, -1.1, -8.1},
  {-2.6, -1.7, -8.4},
  {-2.3, -0.8, -7.5},
  {-0.7, 0.1, -6},
  {0.8, 0.5, -4.4},
  {2.9, 1, -2.5},
  {3.4, 3, 0},
  {3.1, 2.9, 1.3},
  {3.5, 3.8, 2.4},
  {2.7, 4, 1.3},
  {-0.4, 1.5, -2.8},
  {-1.3, 0.2, -4.5},
  {-2.5, 0.1, -5.5},
  {-1.1, 0, -6.6},
  {0, 0.3, -6.8},
  {0.5, 0, -5.3},
  {0.3, 0, -3.9},
  {0, 0, -3.3},
  {0, 0, -2.9},
  {-0.1, 0.2, -2.7},
  {-0.4, 0, -2.8},
  {-0.1, 0.1, -2.8},
  {-0.3, 0.1, -2.5},
  {-0.8, -0.1, -2.7},
  {-1.1, -0.4, -2.9},
  {-1.3, -0.7, -3.9},
  {-1.5, -0.8, -4.5},
  {-1.2, -0.5, -4.2},
  {-0.4, -0.8, -4},
  {1.3, 2.3, -1.3},
  {1.6, 4.1, 1.1},
  {0.4, 3.7, 3.7},
  {0.2, 3.3, 3.3},
  {-0.8, 2, 2.8},
  {-1.6, 0.7, 1.6},
  {-2.1, -0.5, -1.2},
  {-1.8, -0.9, -1.6},
  {-1.9, -0.5, -1},
  {-2.1, -0.5, -0.6},
  {-2.5, -0.8, -0.4},
  {-2.7, -1.7, -1},
  {-2.3, -1.8, -1.2},
  {-2.6, -2.1, -0.9},
  {-2.6, -2.5, -0.8},
  {-2.7, -3, -1.1},
  {-2.9, -3.3, -1},
  {-3, -3.4, -1.1},
  {-3.6, -3.6, -1.3},
  {-4.4, -4.1, -2.3},
  {-5.3, -4, -4.1},
  {-6.2, -3.8, -5.9},
  {-4.7, -3.4, -6.7},
  {-2.1, -2.9, -4.6},
  {-0.7, -1.5, -1.3},
  {-0.2, -0.7, 1},
  {-0.1, 0.8, 2.7},
  {0.9, 0.6, 3.7},
  {0.3, 0.3, 1.5},
  {-2, -0.8, -2},
  {-3.1, -1.3, -4.1},
  {-3.7, -1.8, -6.2},
  {-3.8, -2, -7.2},
  {-3.6, -2.5, -7.9},
  {-3.7, -2.7, -8.8},
  {-4, -2.7, -8.7},
  {-4.1, -2.7, -9.5},
  {-4.5, -2.9, -9.9},
  {-4.6, -3.4, -10},
  {-4.4, -3.8, -10.4},
  {-4.6, -4.1, -11.5},
  {-5, -3.7, -11.6},
  {-4.4, -4.3, -12},
  {-5, -4.2, -12.1},
  {-4.8, -4.2, -12.9},
  {-5, -4.3, -13.1},
  {-2.7, -4, -13.1},
  {0.2, -2.8, -10.3},
  {1.3, -0.5, -6.3},
  {2.9, 0.4, -2.9},
  {4.1, 0.7, -0.2},
  {4.9, 1.2, 1.2},
  {3.9, 1.4, -0.2},
  {-0.5, -0.3, -3.6},
  {-1.1, -1, -6.3},
  {-1.6, -1.3, -7.2},
  {-1.4, -1.3, -7.9},
  {-1.3, -1.3, -9.2},
  {-0.8, -1.8, -9.4},
  {-1.1, -1.7, -9.5},
  {-0.7, -1.8, -10.2},
  {-2.1, -2.1, -10.6},
  {-2.2, -2.3, -11},
  {-2.6, -2.5, -11},
  {-2.5, -2.8, -11.3},
  {-2.4, -2.9, -11.4},
  {-3.1, -3.3, -11.4},
  {-3.3, -3.7, -12.5},
  {-3.7, -3.8, -12.4},
  {-3.9, -4.1, -12.8},
  {-2.1, -3.5, -12.4},
  {1.6, -2.7, -9.7},
  {2.9, -0.4, -6.1},
  {4, 1.6, -2.2},
  {4.3, 2.3, 0.5},
  {4, 2.6, 1.4},
  {4.4, 2.3, 0.2},
  {0.6, 0.2, -3.1},
  {-1.4, -0.4, -5.7},
  {-1.4, -0.7, -6.7},
  {-1.3, -1.1, -8.1},
  {-1.2, -1.2, -8.1},
  {-1.9, -1.5, -9},
  {-2.2, -1.9, -10},
  {-1.8, -2.1, -10.5},
  {-1.6, -2.3, -11.1},
  {-2.1, -2.7, -11.5},
  {-3.1, -3.2, -11.5},
  {-1.9, -3, -11.8},
  {-2.5, -3.4, -12.6},
  {-2.9, -3.4, -12.4},
  {-3.4, -3.2, -13},
  {-2.7, -3.4, -13.1},
  {-3, -3.2, -13.3},
  {-1.2, -2.6, -13.1},
  {1.2, -1.6, -9.9},
  {3.9, 0.7, -5.7},
  {5.1, 1.2, -2.6},
  {4.5, 1.5, -0.1},
  {4.1, 4, 1},
  {2.7, 3.1, 0.2},
  {0, 0.5, -3.3},
  {-1.8, -0.5, -5.2},
  {-2.5, -1.1, -6.9},
  {-3.1, -1.5, -7.7},
  {-3.3, -1.9, -8.6},
  {-3.7, -2.4, -8.9},
  {-3.5, -2.7, -10.1},
  {-4.4, -2.9, -9.9},
  {-4.3, -3.3, -10.9},
  {-4.2, -2.9, -11},
  {-4.5, -3, -11.9},
  {-4.3, -3.4, -12},
  {-3.9, -3.6, -12.6},
  {-4.4, -3.7, -12.4},
  {-4.8, -4.1, -13.1},
  {-5, -4.4, -13.6},
  {-4.8, -4, -13.2},
  {-3.2, -3.5, -13.6},
  {0.1, -2.5, -11.3},
  {2, -0.3, -5.8},
  {2.6, 1.1, -3.4},
  {3, 0.8, -0.4},
  {3.1, 1.6, 1.1},
  {3.4, 2.5, -0.3},
  {-0.4, -0.3, -4.5},
  {-1.9, -1.1, -6.6},
  {-1.9, -1.3, -8.3},
  {-2.3, -1.6, -9},
  {-2.6, -1.8, -9.6},
  {-1.9, -1.9, -10.5},
  {-2.2, -2.1, -10.7},
  {-2.8, -2.3, -11.8},
  {-3.3, -2.7, -11.4},
  {-2.9, -3, -12},
  {-3.1, -2.8, -12.6},
  {-3.7, -3.4, -13.1},
  {-4.1, -3.5, -13.4},
  {-3.8, -4.1, -13.6},
  {-3.6, -4, -13.4},
  {-3.9, -4, -14},
  {-3.6, -3.6, -13.8},
  {-1.8, -3.2, -14.5},
  {0.5, -2.4, -10.4},
  {2.5, 0, -6.5},
  {5.3, 0.5, -3},
  {5.5, 2.7, -0.7},
  {5.4, 2.9, 1},
  {4.6, 2.9, 0.2},
  {0.5, -0.1, -3.7},
  {-1.4, -0.9, -6.3},
  {-1.7, -1.4, -7.6},
  {-2.5, -1.5, -8.8},
  {-2.6, -1.9, -9.7},
  {-1.7, -2.4, -10.5},
  {-3.1, -2.7, -10.6},
  {-3.6, -2.9, -10.6},
  {-4, -3.4, -11.4},
  {-4.2, -3.6, -11.7},
  {-5.3, -4.2, -12.2},
  {-5.2, -4.5, -12.7},
  {-5.3, -4.7, -12.7},
  {-7.3, -5.1, -13.1},
  {-7.2, -5.6, -13.2},
  {-6.9, -5.7, -13.9},
  {-6.9, -5.9, -13.8},
  {-5.1, -5.4, -14.3},
  {-2.9, -5.2, -10.8},
  {-1.6, -2.3, -6.5},
  {-1.3, 0.6, -4.3},
  {-0.7, 0.7, -1.1},
  {-0.3, 0.8, 0},
  {-0.5, 0.3, 0},
  {-3.5, -1.2, -2},
  {-5.4, -2.7, -5.8},
  {-6.5, -3.9, -7.7},
  {-6.9, -4.6, -8.7},
  {-7.2, -5, -9.7},
  {-7.7, -5.4, -10.5},
  {-7.7, -6, -11.1},
  {-7.2, -6.3, -12.3},
  {-7.5, -6.6, -12.6},
  {-8.1, -6.9, -13.2},
  {-7.8, -7.2, -13.1},
  {-7.4, -7.4, -13.7},
  {-7.2, -7.7, -13},
  {-8.1, -7.5, -14.2},
  {-7.9, -7.5, -14.4},
  {-7.8, -8, -14.6},
  {-7.7, -7.9, -14.9},
  {-6.5, -7.1, -14.7},
  {-5.6, -6.3, -11.5},
  {-3.1, -3.8, -6.9},
  {-1, -2, -5},
  {-1.4, -1.7, -2.5},
  {-1.1, -0.5, -1.5},
  {-0.8, -1, -2.2},
  {-3.1, -2.8, -5.2},
  {-5.1, -3.7, -6.7},
  {-6, -4.7, -8.8},
  {-6.1, -5, -9.6},
  {-6.4, -5.7, -10.3},
  {-6.2, -6, -10.7},
  {-5.4, -5.6, -9.8},
  {-4.7, -5.2, -8.7},
  {-4.8, -5.1, -8.1},
  {-5, -5, -7.9},
  {-4.9, -5, -7.7},
  {-5, -4.9, -7.6},
  {-5.3, -5.4, -8.5},
  {-6, -5.5, -9},
  {-5.7, -5.6, -9.5},
  {-5.2, -5.2, -9},
  {-5.1, -5.2, -8.9},
  {-4.9, -3.9, -8},
  {-4.3, -4.2, -6.4},
  {-4.1, -5.1, -4.4},
  {-3.6, -4.7, -2.1},
  {-3.7, -3.7, -0.5},
  {-3.7, -3, 0.1},
  {-3.9, -2.9, -0.5},
  {-3.8, -3.8, -1},
  {-4.3, -3, -1.9},
  {-4.4, -3.2, -3.8},
  {-4.4, -3.2, -3.7},
  {-4.3, -3.7, -3.4},
  {-3.9, -4.2, -3.2},
  {-3.9, -4.5, -3.3},
  {-4, -4.4, -3.2},
  {-4.3, -5.3, -3.4},
  {-3.3, -4.9, -3.9},
  {-2.7, -4.5, -4},
  {-2.1, -4.2, -3.8},
  {-1.8, -3.3, -3.6},
  {-2.1, -2.9, -3.6},
  {-1.6, -2.8, -3.6},
  {-2.8, -2.7, -3.6},
  {-2.9, -2.2, -3.6},
  {-2.7, -1.6, -3.1},
  {-0.9, -1.4, -2.1},
  {1.6, -0.1, -1},
  {3, 0.8, 0.1},
  {4, 2.3, 2.8},
  {3.4, 1.1, 2.5},
  {2.9, 1.2, 1.9},
  {0.2, 2.8, -0.8},
  {-0.2, 2.8, -2.2},
  {0.5, 3, -3.4},
  {0.8, 3.4, -4.2},
  {0.7, 3.4, -5.1},
  {-0.2, 3.3, -5.4},
  {-0.3, 3.4, -5.8},
  {-1.2, 3.3, -6.9},
  {-1.6, 3.1, -7.3},
  {-0.3, 3.1, -7.1},
  {0.5, 3.3, -7.4},
  {0, 3.6, -7.8},
  {-0.7, 3.2, -8.1},
  {-0.9, 3, -8.8},
  {-0.4, 2.6, -9.3},
  {-1.1, 1.5, -9.6},
  {-1.4, 1.6, -10},
  {0.7, 2, -9.6},
  {3.5, 2.6, -6.7},
  {6, 4.9, -3.2},
  {6.4, 7.1, 0},
  {7, 7.4, 2.8},
  {6.7, 8.4, 4.1},
  {6.1, 8.2, 3.2},
  {2.3, 5.2, 0.3},
  {2, 2.7, -2.3},
  {0.1, 1.8, -3.8},
  {-0.4, 1.1, -5.6},
  {-0.8, 0.6, -6.1},
  {-1.1, 0, -7.1},
  {-1.8, 0.3, -6.8},
  {-1.8, 0, -8},
  {-1.4, -0.2, -7.8},
  {-1.6, -0.5, -8.9},
  {-1, -0.6, -8.3},
  {-2.1, -0.6, -9.5},
  {-1.5, -1, -9.3},
  {-1.8, -1, -9.4},
  {-1.8, -1, -10.1},
  {-2, -1.1, -10.1},
  {-1.5, -1.2, -9.9},
  {0.5, -0.8, -10},
  {3, -1, -6.2},
  {4.5, 2.2, -2.7},
  {5.7, 3.4, 0.1},
  {5.4, 5.6, 3.2},
  {5.4, 5.8, 4.4},
  {5, 5.6, 3.7},
  {2.8, 3.2, 0.7},
  {0.8, 0.9, -2.8},
  {0.8, 0.1, -4.1},
  {1.2, -0.4, -5.7},
  {1.5, -0.6, -6.3},
  {0.4, -0.7, -6.7},
  {0, -0.9, -7.4},
  {-1.2, -1.5, -7.8},
  {-0.9, -1.9, -8.3},
  {-0.2, -1.9, -8.7},
  {0, -2, -8},
  {-1.4, -1.7, -8},
  {-0.4, -1.7, -8.7},
  {-0.5, -2.1, -8.4},
  {-1.5, -1.9, -9.1},
  {-1.4, -2.2, -9.9},
  {-1.7, -2.2, -10.2},
  {-1.3, -2.2, -9.4},
  {2.7, -1.2, -6.9},
  {4, 1.5, -3},
  {5.6, 3.1, 0.3},
  {5.4, 4.4, 2.5},
  {4.6, 5.4, 4},
  {4.4, 4.4, 3.2},
  {1.8, 1.9, -0.3},
  {0.2, 0.3, -2.7},
  {-0.5, -0.3, -3.8},
  {-1, -0.7, -4.9},
  {-1.8, -1.2, -6.2},
  {-1.7, -0.3, -7},
  {-1.7, 0.8, -7.3},
  {0, 1.7, -7.7},
  {1.4, 2.3, -8.3},
  {2.3, 1.2, -9.3},
  {0.9, 1.2, -8.4},
  {0.2, 1.2, -9},
  {0.2, 0.9, -9.6},
  {0.3, 1.1, -9.4},
  {0, 1, -10.2},
  {-0.9, 0.7, -10.8},
  {-1, 1.1, -10.8},
  {0.4, 1.2, -10.9},
  {3.4, 2.1, -8.1},
  {3.8, 4.7, -4.3},
  {4.7, 5, -0.6},
  {4.9, 5.3, 2},
  {5, 6.1, 2.7},
  {4.7, 6.3, 4.5},
  {3.1, 5.3, 1.3},
  {1.9, 4.2, -1.4},
  {1.9, 3.6, -3.2},
  {1.5, 3, -4.3},
  {1.1, 3.2, -6.1},
  {0.4, 2.8, -6.2},
  {-0.3, 2.6, -7.3},
  {-0.5, 2.3, -6.8},
  {-0.4, 1.9, -7.3},
  {-0.8, 1.4, -7.7},
  {-0.5, 1.2, -9},
  {-1.3, 1, -9},
  {-2.9, 1, -9.7},
  {-1.3, 0.6, -9.9},
  {-3, 0, -10.3},
  {-4.1, -0.6, -10.4},
  {-3.6, -0.5, -10.3},
  {-0.7, -0.3, -11.2},
  {0.4, 0.2, -7.1},
  {1.1, 2, -3.4},
  {2, 2.8, -0.1},
  {2.4, 3.8, 1.9},
  {0.3, 4.5, 2.7},
  {-0.8, 4.7, 1.4},
  {-3.5, 3.5, -0.2},
  {-4.8, 0.8, -1.2},
  {-5.8, -1.9, -2.5},
  {-6.4, -2.7, -3.7},
  {-7, -3.1, -4.7},
  {-7.7, -3.7, -7.1},
  {-7.6, -4.2, -8.2},
  {-7.4, -4.7, -9.5},
  {-7.1, -5, -9.8},
  {-7.7, -5, -10.4},
  {-7.5, -5.1, -11.8},
  {-7.4, -5.1, -12.3},
  {-7.5, -4.7, -11.9},
  {-7.3, -4.7, -12.5},
  {-8.4, -5.8, -12.9},
  {-8.1, -5.8, -13.3},
  {-7.1, -5.6, -13.7},
  {-4.8, -5.4, -14.2},
  {-2.7, -4.3, -10.8},
  {-1.6, -2.6, -6.6},
  {-1.3, -1.2, -3.7},
  {-0.9, -0.5, -1},
  {-0.9, 0.1, 1.1},
  {-1.8, 0, 0.4},
  {-3.3, -1.5, -1.5},
  {-6.1, -2.8, -5.2},
  {-7, -3.5, -6.7},
  {-6.7, -4.3, -9.2},
  {-6.9, -5.2, -9.9},
  {-7.7, -5.5, -10.7},
  {-7.4, -5.4, -11.5},
  {-7.2, -5.6, -11.9},
  {-6.7, -5.4, -13.1},
  {-7.5, -5.3, -13.1},
  {-7.8, -6.1, -13.6},
  {-8.9, -6.7, -14.3},
  {-9.3, -6.9, -15},
  {-9.2, -6.3, -15},
  {-9.3, -7, -15.7},
  {-9.5, -7.4, -15.9},
  {-8.1, -7.2, -15.8},
  {-5.6, -7.2, -15},
  {-2.2, -6.3, -10.8},
  {-0.7, -3.3, -7.7},
  {-0.2, -2.8, -4.5},
  {-0.4, -2.1, -2.2},
  {-1.8, -2.3, -0.7},
  {-3.1, -2.5, -1.1},
  {-3.4, -3, -2.4},
  {-4.3, -3, -3.7},
  {-4.6, -3.3, -4.5},
  {-5.3, -4, -5.6},
  {-6.1, -4.9, -6.4},
  {-6.2, -4.9, -7.6},
  {-6.2, -5, -7.8},
  {-6.2, -5, -8.5},
  {-6.9, -5.1, -8.6},
  {-6.8, -5.2, -9.3},
  {-8, -5.3, -8.9},
  {-8.4, -6, -9.7},
  {-9.3, -6.4, -11.1},
  {-9.1, -7.2, -11.1},
  {-7.5, -7.6, -12.1},
  {-7.7, -8, -13},
  {-6.2, -7.5, -11.3},
  {-5, -6.7, -9.4},
  {-4.7, -5.2, -7.5},
  {-5.1, -3.7, -6.1},
  {-5.8, -3.1, -4.1},
  {-6.4, -3.1, -3.4},
  {-6.3, -4.1, -2.8},
  {-6.4, -4.9, -3.1},
  {-6.5, -5.3, -3.5},
  {-6.8, -5.5, -3.8},
  {-6.5, -5.5, -3.8},
  {-6.4, -5.6, -3.8},
  {-6.2, -5.3, -3.8},
  {-6.2, -5.1, -3.8},
  {-6, -5.3, -3.8},
  {-4.9, -5.1, -3.8},
  {-4.5, -5, -3.7},
  {-4.5, -5.1, -3.7},
  {-4.3, -5, -3.6},
  {-4.6, -4.7, -3.6},
  {-4.8, -4.8, -3.6},
  {-4.9, -4.7, -3.6},
  {-4.4, -4.6, -3.6},
  {-4.7, -4.6, -3.6},
  {-4.2, -4.1, -3.3},
  {-3.1, -3.4, -2.5},
  {-3.5, -3, -1.9},
  {-3.1, -3.2, -1.6},
  {-2.8, -3.1, -1.5},
  {-3.1, -2.6, -1.4},
  {-2.4, -2.7, -0.6},
  {-1.8, -2.8, -1.1},
  {-1.6, -2.9, -1.5},
  {-2.4, -2.9, -1.6},
  {-2, -2.8, -1.6},
  {-1.1, -2.5, -1.6},
  {-0.9, -2.4, -1.6},
  {-0.9, -2.3, -1.5},
  {-0.9, -1.8, -1.4},
  {-0.8, -1.7, -1.4},
  {-1.1, -1.9, -1.2},
  {-0.8, -1.5, -1.1},
  {-0.6, -1.4, -1.2},
  {-0.3, -1.3, -1.3},
  {-0.2, -1.1, -1.3},
  {-0.5, -1, -1.3},
  {-0.8, -1, -1.2},
  {-0.1, -1, -1.2},
  {0.1, -0.9, -1.2},
  {0.6, -0.3, -0.8},
  {0.9, 0.4, 0.2},
  {1.6, 1, 0.2},
  {1.9, 1.6, 0.7},
  {1.3, 1.9, 1.2},
  {1.6, 1.9, 1.3},
  {2.6, 1.5, 1.2},
  {2.6, 1.2, 0.9},
  {2.8, 0.9, 0.6},
  {3, 1, 0.4},
  {2.8, 1, 0.4},
  {2.7, 0.9, 0.4},
  {2.4, 1, 0.3},
  {2.3, 0.9, 0.2},
  {2.6, 1, 0.2},
  {2.7, 1, -0.6},
  {2.6, 1.1, -1},
  {3, 1, -1.1},
  {2.9, 0.7, -0.8},
  {3.1, 0.8, -0.6},
  {2.8, 1.1, -0.4},
  {3, 0.9, -0.4},
  {2.7, 1.1, -0.6},
  {1.8, 1.3, -0.7},
  {2.6, 1.8, -0.5},
  {2.9, 2.3, 0.3},
  {3.5, 3.1, 0.9},
  {3.4, 3.6, 1.4},
  {3.8, 3.7, 2},
  {4.3, 3.8, 2.1},
  {3.8, 3.8, 2.4},
  {3.1, 3.3, 1.7},
  {2.9, 2.5, 1.6},
  {3.7, 2.1, 0.9},
  {3.2, 2, 0.6},
  {3.1, 1.9, 0.5},
  {2.9, 1.9, 0.3},
  {3, 1.9, 0.1},
  {3, 2, 0.1},
  {3.1, 1.8, -0.4},
  {3.1, 1.8, 0},
  {3.1, 2.1, 0},
  {3.1, 2.2, 0.1},
  {2.8, 2.4, 0},
  {3, 2, -0.1},
  {2.4, 1, -0.3},
  {1.7, 0.8, -0.2},
  {1.4, 1, 0},
  {2.3, 1, 0.4},
  {3.6, 2.3, 0.6},
  {4.5, 5.1, 0.9},
  {6, 5.6, 1.6},
  {7.9, 6.1, 3},
  {7.9, 7, 5.6},
  {7.3, 6.6, _},
  {5.8, 5.3, _},
  {4.2, 3.5, _},
  {3.3, 3.3, _},
  {2.6, 3, _},
  {3.2, 2.8, _},
  {2.9, 2.7, _},
  {2.5, 2.5, _},
  {1.7, 1.9, _},
  {2.1, 1.7, _},
  {1.2, 1.5, _},
  {1.5, 1.1, _},
  {0.9, 1.5, _},
  {0.7, 0.8, _},
  {0.5, 0.7, _},
  {0.9, 1.1, _},
  {0.2, 0.9, _},
  {0.6, 0.9, _},
  {3.3, 1.9, _},
  {5.4, 2.9, _},
  {7.4, 5, _},
  {8.4, 6.1, _},
  {8.4, 6.8, _},
  {9, 6.9, _},
  {8.2, 7.4, _},
  {6.5, 6.3, _},
  {5.1, 4.6, _},
  {3.9, 3.6, _},
  {3.6, 3.3, _},
  {3.5, 3.2, _},
  {3.1, 3.5, _},
  {3.7, 2.9, _},
  {3.6, 3, _},
  {3.5, 2.9, _},
  {3.3, 2.2, _},
  {2.2, 2.1, _},
  {2, 2, _},
  {3, 1.6, _},
  {2, 1.4, _},
  {2.2, 0.9, _},
  {1.9, 1.1, _},
  {3.2, 1.5, _},
  {6, 2.4, _},
  {6.6, 3.9, _},
  {7.6, 6.2, _},
  {10, 7.8, _},
  {11.6, 7.9, _},
  {11.2, 8.6, _},
  {8.1, 8.8, _},
  {6.7, 6.9, _},
  {6.1, 5, _},
  {5.7, 4.2, _},
  {5.2, 3.8, _},
  {4.8, 3.6, _},
  {4.5, 3.9, _},
  {3.6, 3.1, _},
  {3, 3.2, _},
  {3.2, 3.4, _},
  {2.5, 2.6, _},
  {2.3, 2.5, _},
  {2.4, 1.7, _},
  {1.9, 1.7, _},
  {1.2, 1.2, _},
  {1.3, 1.3, _},
  {1.5, 0.7, _},
  {2.3, 0.8, _},
  {4.8, 1.7, _},
  {6.6, 2.4, _},
  {8.7, 4.9, _},
  {11.1, 7.2, _},
  {11.1, 9.6, _},
  {11, 10.2, _},
  {9, 9.8, _},
  {5.9, 7.5, _},
  {4.1, 5.1, _},
  {3, 3.8, _},
  {2.5, 3.1, _},
  {2.1, 2.9, _},
  {2.3, 3.4, _},
  {2.9, 3.2, _},
  {2.8, 3.1, _},
  {2, 2.2, _},
  {1.5, 1.8, _},
  {0.2, 1.5, _},
  {0.2, 1.1, _},
  {0.3, 0.9, _},
  {-0.1, 0.7, _},
  {-0.2, 0.6, _},
  {0.3, 0.3, _},
  {-0.4, 0.4, _},
  {3.3, 0.8, _},
  {5.6, 2.2, _},
  {6.8, 4.2, _},
  {7.8, 5.4, _},
  {7.2, 7.1, _},
  {8, 9.1, _},
  {7.8, 8.7, _},
  {3.8, 7.3, _},
  {1.8, 4.1, _},
  {1.5, 2.7, _},
  {0.7, 2.1, _},
  {0, 1.4, _},
  {-0.3, 1.3, _},
  {0, 1, _},
  {-0.1, 1, _},
  {0.4, 1, _},
  {0.3, 0.7, _},
  {0.1, 0, _},
  {-0.7, -0.1, _},
  {-1.3, -0.6, _},
  {-1.8, -0.7, _},
  {-2.2, -0.7, _},
  {-2.4, -1.1, _},
  {-1.3, -0.9, _},
  {1.5, -0.3, _},
  {3.7, 0.8, _},
  {5.3, 2.8, _},
  {5.9, 3.6, _},
  {5.4, 5.1, _},
  {5.5, 7.3, _},
  {6.1, 7.7, _},
  {3, 6.1, _},
  {0.4, 2.9, _},
  {-0.3, 1.5, _},
  {-0.7, 0.9, _},
  {-0.8, 0.3, _},
  {-0.8, 0.3, _},
  {-1.1, 0.1, _},
  {-1, -0.3, _},
  {-1.3, -0.5, _},
  {-1.9, 0, _},
  {-2.2, -0.2, _},
  {-2.7, -0.9, _},
  {-2.7, -1.1, _},
  {-3.9, -1.3, _},
  {-2.3, -1.9, _},
  {-3.5, -1.9, _},
  {-3.3, -2.2, _},
  {-1, -1.8, _},
  {0, -0.9, _},
  {-0.8, 1.8, _},
  {0, 1.9, _},
  {0.2, 2.1, _},
  {-0.2, 2.6, _},
  {-1.1, 1.6, _},
  {-2.1, 0.6, _},
  {-3.3, -0.5, _},
  {-4.3, -1, _},
  {-4.7, -1.6, _},
  {-4.8, -2.2, _},
  {-4.7, -2.6, _},
  {-4.5, -2.9, _},
  {-4.5, -3, _},
  {-4.7, -3.3, _},
  {-4.7, -2.9, _},
  {-4.9, -2.7, _},
  {-5, -2.9, _},
  {-5, -3.5, _},
  {-5, -3.4, _},
  {-5.4, -3.7, _},
  {-5.3, -3.9, _},
  {-5.1, -3.5, _},
  {-5, -2.9, _},
  {-4.8, -2.2, _},
  {-3.8, -1.2, _},
  {-3.2, -0.4, _},
  {-2.9, 0.4, _},
  {-2.6, 0.8, _},
  {-2.9, 0.4, _},
  {-3.8, -0.6, _},
  {-4.9, -1.8, _},
  {-5.9, -2.5, _},
  {-6.5, -2.7, _},
  {-7, -2.9, _},
  {-7.5, -3.4, _},
  {-7.6, -4.1, _},
  {-7.7, -4.4, _},
  {-7.6, -4.4, _},
  {-7, -4.2, _},
  {-7, -4.5, _},
  {-6.5, -5.2, _},
  {-6.7, -5.6, _},
  {-7.1, -5.8, _},
  {-7.6, -6.1, _},
  {-7.2, -6.3, _},
  {-6.8, -6.1, _},
  {-4.1, -5.3, _},
  {-2.6, -3.6, _},
  {-2.4, -2, _},
  {-1.5, -1, _},
  {-0.8, 0, _},
  {-0.2, 0.7, _},
  {0, 1.1, _},
  {-1.3, 0.5, _},
  {-3.1, -1.2, _},
  {-3.8, -1.8, _},
  {-4.1, -2.1, _},
  {-4.2, -2.6, _},
  {-4.1, -2.9, _},
  {-3.8, -3.1, _},
  {-2.7, -3.4, _},
  {-2.2, -3.3, _},
  {-1.5, -3.2, _},
  {-1.8, -3.3, _},
  {-1.8, -3.1, _},
  {-1.7, -2.8, _},
  {-2.3, -3.4, _},
  {-1.7, -3.5, _},
  {-2.3, -3.5, _},
  {-1.9, -2.9, _},
  {-0.5, -1.8, _},
  {0.4, -1, _},
  {0.8, -0.7, _},
  {1.6, 0.2, _},
  {0.9, 1.6, _},
  {0.4, 1.7, _},
  {-0.6, -0.1, _},
  {-0.9, -0.5, _},
  {-0.7, -0.9, _},
  {-1.7, -1.1, _},
  {-1.4, -1.3, _},
  {-1.3, -1.9, _},
  {-2.7, -2, _},
  {-2.6, -2.2, _},
  {-2.5, -2.6, _},
  {-2.4, -2.5, _},
  {-2.5, -2.3, _},
  {-3, -2.3, _},
  {-3.7, -2.5, _},
  {-3.9, -2.3, _},
  {-3.1, -2.5, _},
  {-2.5, -1.9, _},
  {-3, -2.3, _},
  {-1.8, -2.6, _},
  {1.1, -2.2, _},
  {3.3, -0.2, -4},
  {3.9, 3, -2.8},
  {4.4, 6.1, 0.2},
  {4.8, 6.1, 3.6},
  {4.6, 6.5, 5.2},
  {4.4, 5.6, 6.5},
  {2.8, 3.5, 4.3},
  {-0.6, 2.1, 1.2},
  {-1.8, 1.1, -1.7},
  {-1.6, 0.3, -2.9},
  {-1.3, 0.1, -3.9},
  {-1.1, 0.3, -4.4},
  {-1.8, 1, -4.5},
  {-2, 1.2, -4.6},
  {-0.9, 1.1, -5.7},
  {-1.3, 0.1, -7.3},
  {-2.8, -0.2, -8.6},
  {-3, -0.7, -9.3},
  {-3.3, -1.2, -10.1},
  {-3.3, -1.5, -10.7},
  {-3.3, -1.9, -11.3},
  {-2.9, -2, -12.3},
  {-2.9, -1.8, -12.4},
  {-0.5, -1, -12},
  {1.5, 0.3, -6.8},
  {2, 1.9, -3.1},
  {2.5, 2.9, 1},
  {2.9, 3.5, 4.4},
  {3.4, 4.1, 6.1},
  {3.3, 4.6, 5.3},
  {1.7, 4.1, 2.8},
  {-1.2, 2, -1.4},
  {-2.2, 1.2, -4.1},
  {-2.6, 0.9, -6},
  {-2.6, 0.3, -6.8},
  {-3, 0, -8},
  {-3.5, -0.8, -8.6},
  {-3.6, -1.5, -9.7},
  {-4.1, -1.9, -10.2},
  {-4.1, -2, -11.1},
  {-3.6, -2.1, -11.3},
  {-4.4, -1.9, -11.8},
  {-3.7, -2, -12.7},
  {-3.7, -2.2, -12.8},
  {-4.3, -2.8, -13},
  {-4.4, -2.7, -14.4},
  {-3.9, -2.4, -13.8},
  {-1, -1.3, -12.7},
  {0.6, 0, -8.2},
  {1.4, 2, -2.8},
  {2.1, 3, 0.3},
  {2.3, 3.6, 3.5},
  {2.9, 4.8, 7.1},
  {2.8, 5, 5.6},
  {1.3, 4.1, 1.8},
  {-0.8, 1.3, -1.4},
  {-0.5, 0.4, -4.2},
  {-1.3, 0.1, -6.1},
  {-1.9, -0.5, -8.1},
  {-3.9, -1, -8.6},
  {-4.5, -1.6, -9.6},
  {-4.5, -1.9, -10.2},
  {-4.8, -2.2, -10.6},
  {-4.8, -3, -11.5},
  {-5.1, -3.4, -11.5},
  {-6.4, -4.1, -12.1},
  {-6.2, -4.7, -12.2},
  {-7, -5, -13.5},
  {-7.1, -5.5, -13.1},
  {-7.3, -5.7, -14.4},
  {-7.2, -5.6, -14.4},
  {-3.1, -4.7, -13.7},
  {-1.4, -2.8, -7.8},
  {-0.5, -1.2, -4.3},
  {1.4, 0.6, -0.4},
  {1.9, 1.7, 2.3},
  {1.4, 2.6, 5.3},
  {1.8, 3.8, 5},
  {-0.1, 2.4, 2.9},
  {-1.6, 0.6, 0.8},
  {-3.2, -0.4, -3.2},
  {-3.7, -0.9, -5.3},
  {-4.5, -1.5, -6.2},
  {-5, -2.3, -7.7},
  {-5.1, -2.9, -9},
  {-5.8, -3.2, -9.3},
  {-5.7, -3.3, -10.4},
  {-6.3, -3.8, -11.3},
  {-6.5, -3.9, -11.6},
  {-6.5, -4, -12},
  {-6.8, -4.7, -12.6},
  {-6.7, -5.1, -13},
  {-7.1, -5.3, -14.3},
  {-7.2, -5.9, -14.2},
  {-6.4, -4.6, -13.8},
  {-2.1, -4.5, -12.7},
  {-0.5, -3.2, -7.8},
  {0.8, -0.3, -4.3},
  {1.1, 0.8, 0.1},
  {1.4, 2.2, 2.5},
  {2.3, 3.6, 4.8},
  {1.9, 4, 4.8},
  {0.2, 2.7, 3.2},
  {-2, 0.3, -1.5},
  {-3.1, -0.7, -4.3},
  {-3.4, -1.1, -5.7},
  {-3.6, -1.4, -6.8},
  {-4.1, -2, -8.3},
  {-4.8, -2.3, -9},
  {-4.5, -2.4, -8.6},
  {-4.9, -3, -9.5},
  {-5.5, -3.5, -10.5},
  {-6.1, -3.9, -11.2},
  {-6.1, -4.2, -11.7},
  {-6.3, -4.3, -12.3},
  {-6.5, -4.7, -12.3},
  {-6.7, -4.7, -12.6},
  {-6.4, -4.6, -13.6},
  {-5.7, -4.7, -14.1},
  {-1.8, -4.3, -12.7},
  {0.5, -2.3, -7.6},
  {1.4, 0.9, -3.2},
  {1.8, 2.1, 0.6},
  {3.1, 3.5, 3.6},
  {3.1, 4.4, 4.8},
  {3, 4.5, 5.3},
  {1.2, 3, 3.4},
  {-0.5, 0.9, 0.4},
  {-0.7, 0.3, -2.4},
  {-0.9, -0.2, -3.8},
  {-2.2, -0.4, -5.1},
  {-1.5, -0.7, -6.2},
  {-1.6, -1, -6.3},
  {-1.6, -1.2, -7.3},
  {-2, -1.5, -8.2},
  {-1.4, -2, -8.2},
  {-2.1, -2.4, -8.5},
  {-2.3, -2.7, -8.1},
  {-2.5, -2.6, -6.9},
  {-2.9, -2.6, -8},
  {-2.5, -2.4, -8.1},
  {-2.9, -2.6, -8.4},
  {-1.7, -2.2, -8.7},
  {-0.5, -1.6, -7.1},
  {-0.4, -1.2, -3.7},
  {-0.9, -1, -1.3},
  {-0.6, -0.1, -0.4},
  {-0.1, 0.2, 0.1},
  {-0.8, 0, 1.6},
  {-1.1, -0.1, 2.1},
  {-0.4, -0.7, 1.7},
  {-0.2, -0.7, 0.6},
  {-0.2, -0.8, 0},
  {-0.8, -1.3, 0},
  {-0.3, -1.3, -0.3},
  {0, -1.2, -0.8},
  {-0.8, -1.3, -0.4},
  {-0.9, -1.5, -0.6},
  {-1.2, -1.4, -0.6},
  {-0.3, -1.5, -1},
  {-0.7, -1.7, -1.2},
  {-0.6, -1.8, -1.2},
  {-0.1, -1.5, -1},
  {0.1, -1.8, -1},
  {1.1, -1.7, -1.4},
  {0, -1.7, -1.1},
  {-0.7, -1.5, -0.9},
  {1, -1.4, -0.1},
  {2.3, -1, 0.9},
  {3.1, -0.8, 2.2},
  {3.1, -0.5, 2.9},
  {3.4, 0, 3.1},
  {3.9, 0.1, 3.7},
  {2.2, 1, 4.2},
  {0.4, 0.5, 3.4},
  {0.8, 0.3, 2.6},
  {0.6, 0.6, 1.9},
  {1.1, 0.8, 1.6},
  {2.4, 0.9, 1.3},
  {2.4, 0.9, 1.2},
  {2.1, 0.9, 1.2},
  {2, 0.7, 1},
  {2.3, 0.6, 0.9},
  {2.2, 0.6, 0.5},
  {2.7, 0.2, 0.1},
  {2.5, 0, -0.2},
  {2, -0.1, -0.3},
  {0.5, -0.2, -0.1},
  {0.7, 0.2, 0.3},
  {0.4, 0.6, 0.6},
  {0.4, 0.2, 0.9},
  {0.7, 0.9, 1.7},
  {0.7, 1.8, 2.6},
  {2.3, 1.6, 3.5},
  {5.4, 4.2, 4.8},
  {6.5, 6.4, 6.9},
  {7.4, 8.1, 8},
  {5, 8.1, 6.9},
  {5, 6.6, 5.1},
  {4.4, 4.6, 5.1},
  {2.7, 4, 3.1},
  {2.9, 3.5, 1.7},
  {3.3, 2.5, 0.4},
  {2.8, 1.8, -0.6},
  {1.2, 1.4, -2.2},
  {0, 0.8, -3},
  {0.2, 0.6, -3},
  {-0.3, 0.4, -3.6},
  {0.2, 0, -3.8},
  {0.8, -0.1, -4.4},
  {0.5, -0.3, -5},
  {3.1, -0.4, -4.6},
  {3.3, -0.4, -4},
  {2.6, -0.3, -3.1},
  {2.1, 0, -2},
  {2.6, 0.3, -1.3},
  {2.4, 0.6, -0.5},
  {2.7, 0.5, 0.4},
  {2.5, 1.1, 0.9},
  {2, 1.3, 1.2},
  {2, 1.2, 0.9},
  {2, 0.6, 1},
  {1.6, 1, 0.7},
  {0.5, 0.4, 0.2},
  {0.2, 0.3, 0.1},
  {0.6, 0.3, 0.3},
  {1.5, 0.3, 0.2},
  {1.6, 0.4, 0.1},
  {1.3, 0.4, 0.1},
  {0.4, 0.3, 0},
  {-0.4, 0.4, -0.1},
  {-0.7, 0, 0},
  {-1.1, 0.1, 0.1},
  {-1, -0.1, 0},
  {-1.1, -0.1, -0.2},
  {-1, -0.1, -0.2},
  {-0.9, -0.1, -0.4},
  {-1, -0.2, -0.6},
  {-0.8, 0, -0.6},
  {0.5, 0.5, -0.5},
  {0.5, 0.5, -0.4},
  {1.1, 1, -0.1},
  {1.3, 0.7, 0},
  {1.7, 0.4, 0.2},
  {2.1, 0.3, 0.3},
  {3, 0.5, 0.3},
  {3, 1, 0.3},
  {2.9, 1, 0.1},
  {3, 1, 0.1},
  {3.2, 1, 0.1},
  {3, 1, 0.1},
  {3.4, 1.1, 0.1},
  {3.1, 1.1, 0.1},
  {3.1, 1.4, 0.1},
  {2, 1.4, 0.1},
  {1.6, 1.2, 0.2},
  {1.2, 0.7, 0.2},
  {1.7, 0.6, 0.1},
  {1.2, 0.7, 0},
  {1.4, 1.4, 0.1},
  {1.4, 1, 0.1},
  {1.8, 1.4, 0.1},
  {2.4, 1.6, 0.2},
  {2.4, 1.5, 0.4},
  {2.5, 1.6, 0.8},
  {2.7, 1.7, 0.8},
  {2.3, 2.2, 1},
  {2.1, 1.9, 1.1},
  {1.5, 2, 1.5},
  {1.3, 2.1, 1.4},
  {1.4, 2, 1.6},
  {1.5, 1.7, 1.2},
  {1.5, 1.6, 0.9},
  {1.2, 1.6, 0.8},
  {1.4, 1.7, 0.7},
  {1.3, 1.6, 0.6},
  {1.1, 1.5, 0.4},
  {0.6, 1.3, 0.4},
  {0.4, 1, 0.3},
  {0.4, 1.2, 0.4},
  {0, 1.2, 0.2},
  {0.1, 1.2, 0.2},
  {0.4, 1.2, 0.2},
  {0.4, 1.1, 0.1},
  {0.4, 1, 0.2},
  {0.6, 1, 0.1},
  {1, 1.6, 0.4},
  {1.9, 1.8, 0.7},
  {1.8, 2.2, 1.2},
  {2.2, 2.4, 1.9},
  {1.8, 2.7, 2.1},
  {0.9, 3.3, 2.5},
  {0.8, 3.8, 2.8},
  {1.5, 3.3, 2.5},
  {1.5, 2.7, 2.3},
  {1.3, 2, 2.1},
  {1.4, 1.6, 1.6},
  {1.4, 1.7, 1.2},
  {1, 1.7, 1},
  {1.6, 1.7, 0.8},
  {1.8, 1.4, 0.8},
  {1.8, 1.8, 0.5},
  {1.7, 1.9, 0.6},
  {1.5, 1.9, 0.5},
  {1.3, 1.7, 0.4},
  {1.2, 1.8, 0.4},
  {0.8, 1.7, 0.4},
  {0.4, 1.7, 0.4},
  {0.6, 1.6, 0.5},
  {0.5, 1.6, 0.3},
  {1.2, 1.5, 0.5},
  {1.2, 1.9, 0.7},
  {1.9, 2.4, 1.2},
  {1.9, 3.1, 2},
  {1.4, 3.5, 2.4},
  {1.1, 3.9, 3.3},
  {1.5, 4.2, 3.1},
  {1.6, 3.6, 2.5},
  {1.5, 2.9, 2.4},
  {1.1, 2.4, 1.9},
  {1, 1.9, 1.5},
  {0.9, 1.3, 1.1},
  {0.9, 1.5, 0.9},
  {0.8, 1.3, 0.9},
  {0.7, 1.3, 0.9},
  {0.7, 1.6, 0.7},
  {0.8, 1.1, 0.7},
  {0.8, 1.4, 0.7},
  {0.6, 1.5, 0.6},
  {0.6, 1.2, 0.6},
  {0.4, 0.9, 0.5},
  {0.7, 1, 0.5},
  {0.4, 0.9, 0.6},
  {-0.4, 0.9, 0.5},
  {-0.1, 1.3, 0.8},
  {1.1, 1.5, 0.8},
  {2.4, 3, 1.3},
  {3.1, 4.1, 2.8},
  {3.2, 4.9, 3.8},
  {3.7, 4.8, 5.2},
  {4.5, 5.4, 5.8},
  {4.9, 5.7, 7},
  {4.2, 5, 6.4},
  {2.4, 3.5, 4.8},
  {1.1, 2.7, 3.1},
  {1.6, 1.7, 1.6},
  {1.5, 1.6, 0.6},
  {1.1, 1.9, -0.1},
  {0.8, 1.4, -0.2},
  {0.7, 0.9, -0.4},
  {0.7, 1, -1.2},
  {0.8, 0.9, -1.5},
  {1.1, 0.8, -1.7},
  {1.2, 1, -1.5},
  {1.2, 0.9, -0.9},
  {1, 0.8, -0.6},
  {0.7, 1, -0.5},
  {0.5, 1.1, -0.4},
  {-0.1, 1.7, -0.2},
  {0.1, 2.1, 0},
  {-0.9, 2.9, 0.6},
  {0.3, 2.6, 1.2},
  {0.9, 2.9, 2},
  {0.9, 2.6, 2},
  {1.8, 3.2, 2.6},
  {2.2, 3.5, 2.3},
  {1.8, 3.3, 2.3},
  {0.9, 2.5, 1.8},
  {0.6, 2.5, 1.3},
  {0.7, 2.4, 1.2},
  {1.5, 2.4, 1.1},
  {1.4, 2.4, 1},
  {1.1, 2.4, 0.9},
  {0.6, 2.5, 0.8},
  {0.4, 2.4, 0.6},
  {0.5, 2.2, 0.7},
  {0.8, 2.3, 0.7},
  {1, 2.3, 0.6},
  {0.8, 2, 0.6},
  {0.7, 1.8, 0.5},
  {0.3, 1.7, 0.7},
  {0, 1.7, 0.5},
  {0.2, 2.2, 0.7},
  {0.2, 2.3, 1.1},
  {0.3, 2.6, 1.8},
  {0.5, 2.4, 2.5},
  {0.6, 2.4, 3.1},
  {0.6, 2.3, 2.7},
  {0.6, 2.1, 2.6},
  {0.2, 1.4, 2.5},
  {0.1, 1.2, 2.4},
  {0.1, 0.9, 2.4},
  {0, 0.9, 2.2},
  {-0.4, 0.8, 1.6},
  {-0.7, 0.7, 1.2},
  {-0.7, 0.7, 0.9},
  {-0.5, 0.6, 0.8},
  {-0.6, 0.5, 0.7},
  {-1, 0.4, 0.6},
  {-0.9, 0.3, 0.5},
  {-0.9, 0.4, 0.5},
  {-1.2, 0.4, 0.4},
  {-1.3, 0.4, 0.3},
  {-1.2, 0.3, 0.2},
  {-1.3, -0.1, 0.2},
  {-1.2, -0.1, 0.3},
  {-1.1, 0.5, 0.6},
  {-0.9, 0.8, 1.2},
  {-0.8, 1.3, 2},
  {-0.1, 1.4, 2.7},
  {-0.2, 1.9, 3.9},
  {0.2, 2.3, 4},
  {0.6, 2.4, 3.6},
  {0.5, 2.3, 3.9},
  {0.3, 2.1, 3.6},
  {0.3, 1.7, 2.6},
  {0.3, 1.3, 2},
  {0, 1, 1.6},
  {0, 1.2, 1.3},
  {0, 0.9, 1.2},
  {0, 0.6, 1},
  {0, 0.2, 0.8},
  {0, 0.2, 0.6},
  {-0.1, 0.3, 0},
  {-0.2, 0.4, -0.1},
  {-0.4, 0.4, -0.1},
  {-0.7, 0.1, 0},
  {-1.4, -0.4, -0.1},
  {-1.2, -0.9, -0.3},
  {-1.6, -1.3, -0.3},
  {-1.5, -1.2, 0.1},
  {-0.3, -0.8, 0.6},
  {0.5, 0.4, 1.8},
  {1.3, 1.7, 4},
  {2.1, 2.8, 5.4},
  {2.3, 3.5, 6.4},
  {2.6, 4.1, 6.5},
  {2.6, 4.6, 5.7},
  {1.6, 4.9, 5.7},
  {-0.1, 2.9, 3.6},
  {-1.1, 1.3, 2.1},
  {-1.8, 0.2, 0.1},
  {-2, 0.1, -0.1},
  {-2.3, 0.2, 0.4},
  {-2, -0.2, 0.7},
  {-2.3, -1, 1.3},
  {-2.4, -1.6, 1},
  {-2.9, -2.1, 0.6},
  {-3.1, -2.7, 0.2},
  {-3.2, -3.3, 0.1},
  {-3.6, -3.9, 0},
  {-4.1, -4.3, -0.4},
  {-4.7, -4.7, -0.8},
  {-4.9, -4.9, -0.9},
  {-4.7, -4.3, -0.9},
  {-4.8, -3.8, -0.8},
  {-4.6, -2, -0.1},
  {-4.1, -0.4, 0.7},
  {-3.1, 0.7, 1.3},
  {-3.2, 0.6, 1.1},
  {-3, 0, 0.6},
  {-2.3, -0.1, 0.8},
  {-3, -0.3, 0.9},
  {-3.3, -0.8, 0.7},
  {-3.6, -1, 0.4},
  {-4, -1.6, 0.2},
  {-4.3, -1.9, 0},
  {-4.6, -2.3, -1.1},
  {-5.8, -3, -2.3},
  {-4.8, -3.1, -3},
  {-4.2, -2.7, -2.2},
  {-4, -2.2, -1.7},
  {-4, -2.4, -1.6},
  {-4.1, -2.6, -1.7},
  {-4.2, -2.8, -1.7},
  {-4.3, -2.8, -1.7},
  {-4.3, -2.9, -1.5},
  {-4.5, -3, -1.6},
  {-3.9, -2.7, -2},
  {-3.7, -2.4, -1.8},
  {-2.5, -1.3, -0.7},
  {-0.9, -0.4, 0.3},
  {-0.4, 0.9, 1.3},
  {0.2, 2, 3},
  {0.1, 2.2, 2.8},
  {-0.8, 1.4, 2.2},
  {-1.1, 0.6, 1},
  {-1.8, -0.1, -0.2},
  {-2.4, -0.7, -1.6},
  {-2.5, -1.2, -2.7},
  {-2.6, -1.1, -3.2},
  {-3.3, -0.9, -3.2},
  {-4.1, -1, -3.5},
  {-4.2, -1.8, -4.1},
  {-3.9, -2.7, -3.3},
  {-3.9, -3.1, -2.7},
  {-4.3, -3, -3.3},
  {-4.3, -3.2, -3.4},
  {-4.6, -3.8, -2.7},
  {-4.8, -3.8, -2.4},
  {-5, -3.7, -1.9},
  {-5.1, -3.9, -2.3},
  {-5.1, -4.2, -3.1},
  {-3.9, -3.7, -1.7},
  {-2.7, -2, 0.2},
  {-0.8, -0.7, 1.7},
  {0, 1.5, 4.1},
  {0.1, 2.2, 4.1},
  {-0.7, 1.9, 3.5},
  {-1.5, 3.2, 2.8},
  {-1.4, 2.3, 1.9},
  {-1.9, 0.6, 2.3},
  {-2.7, 0.1, 1.9},
  {-3.7, -0.3, -0.9},
  {-4.6, -0.9, -2.4},
  {-4.5, -1.2, -3},
  {-5, -1.7, -4.4},
  {-5.2, -2.9, -5.3},
  {-5.2, -3.5, -5.8},
  {-4.7, -3.5, -5.4},
  {-4.3, -3.5, -5.2},
  {-3.6, -3.6, -5.1},
  {-3.2, -4, -5.9},
  {-4.2, -4.7, -5.2},
  {-4.5, -5.2, -6.1},
  {-2.9, -4.6, -5.8},
  {-2, -4.1, -4.5},
  {-1.6, -2.6, -3},
  {-0.8, -0.3, -1.5},
  {0, 0.9, 1.5},
  {2.1, 2.2, 2.9},
  {3, 3.8, 5.3},
  {3.6, 4.9, 6.3},
  {3.6, 5.2, 5},
  {3.7, 4.6, 4},
  {2.5, 2.4, 3.1},
  {2.4, 1.1, 1.9},
  {1.8, 0.6, -0.2},
  {2, 1.1, -1},
  {1.8, 1.1, -0.7},
  {1.8, 1.2, -0.1},
  {1.8, 1.3, 0},
  {1.8, 1.1, 0},
  {2, 0.5, 0},
  {1.9, 0.3, 0},
  {0.7, 1.3, -0.2},
  {1.7, 1.5, -0.2},
  {2.8, 1.7, -0.2},
  {2.9, 2, -0.2},
  {2.9, 2.8, 0},
  {3.4, 2.7, 0.4},
  {3.7, 3.6, 1.4},
  {4.3, 3.5, 2.1},
  {4.7, 4.2, 2.7},
  {5.3, 4.1, 3.5},
  {5.9, 5, 5.3},
  {6.7, 7.1, 7},
  {6.8, 7.9, 8.8},
  {6.6, 8.3, 8.1},
  {6.5, 7.7, 7.9},
  {6.4, 7.9, 7.9},
  {6.5, 8, 5.8},
  {6.6, 7.7, 4.3},
  {6.5, 7.2, 3.8},
  {6.2, 7.6, 3.4},
  {6.5, 7.8, 3.4},
  {6.5, 7.8, 3.7},
  {6.7, 8, 4.6},
  {6.2, 7.9, 4},
  {5.5, 7.6, 3.2},
  {5.1, 6.5, 2.8},
  {4.6, 5.1, 2.4},
  {4.7, 4.4, 2.5},
  {4.5, 4.1, 2.4},
  {4.4, 4.2, 2.4},
  {3.6, 4.2, 2.5},
  {3, 3.3, 2.6},
  {3.5, 1.3, 2.6},
  {3.4, 1.3, 2.9},
  {2.9, 2.2, 3.7},
  {2.6, 3.4, 4.8},
  {2.5, 4, 6.3},
  {2.6, 3.6, 6.7},
  {1.8, 2.7, 6.5},
  {0.9, 2, 5.9},
  {0.5, 1.5, 5.6},
  {0.5, 1.3, 4.9},
  {-0.1, 0.9, 4.4},
  {-0.7, 0.4, 4},
  {-0.8, -0.1, 3.5},
  {-2.3, -0.6, 3},
  {-3.1, -1.1, 2.1},
  {-4.1, -1.3, 0.4},
  {-4.9, -1.5, -1.3},
  {-5, -1.7, -3.3},
  {-5.4, -2.2, -4.6},
  {-5.7, -2.5, -5.3},
  {-5.3, -2.7, -5.7},
  {-2.2, -2.6, -5.6},
  {-0.9, -0.8, -2.1},
  {0.4, 1.3, 0.5},
  {1.4, 2.5, 3.2},
  {2.3, 3.4, 3.9},
  {2.7, 4.1, 5.9},
  {2.8, 4.3, 6.5},
  {2.8, 4.3, 7},
  {2.1, 3.5, 6.5},
  {0.7, 2.2, 5.5},
  {-0.1, 1, 4.5},
  {-1.1, 0.6, 3.7},
  {-1.4, -0.2, 2.2},
  {-1.5, -0.8, 0.2},
  {-2.9, -1.3, -1.2},
  {-4.1, -2.3, -3.1},
  {-4.8, -2.6, -4.4},
  {-5.3, -3.2, -5.5},
  {-5.1, -3.5, -6.3},
  {-5.3, -3.8, -6.3},
  {-6, -4, -5.5},
  {-6.3, -4.3, -6.2},
  {-6.5, -3.7, -6.7},
  {-5.7, -3.4, -7},
  {-3, -1.8, -6.9},
  {-0.5, -0.4, -3.5},
  {0.9, 1.6, 0.1},
  {1.8, 2.6, 3.1},
  {2.2, 3.4, 5.2},
  {2.6, 4.2, 5.6},
  {2.5, 4.2, 5.4},
  {2.3, 4, 5.6},
  {1.7, 3.8, 5.7},
  {0.4, 2.4, 4.7},
  {-1.1, 0.8, 2.4},
  {-1.4, 0, 0},
  {-2.4, -1, -1.4},
  {-3.1, -1.6, -1.8},
  {-3.3, -1.9, -3.5},
  {-4.4, -2.4, -4.6},
  {-4.9, -3, -5.4},
  {-5.2, -3.8, -6.8},
  {-5.4, -4.2, -7.3},
  {-6.2, -4.9, -8.2},
  {-6.5, -5.3, -8.2},
  {-5.9, -5.2, -7.8},
  {-6.5, -5.3, -7.9},
  {-6.6, -5.7, -8.3},
  {-4.2, -5.1, -8.1},
  {-1.5, -3.6, -4.5},
  {-0.4, -1, -1.4},
  {0.4, 0, 1.8},
  {1, 1.8, 3.2},
  {1.2, 2.5, 4.6},
  {1.6, 3.5, 4.7},
  {1.6, 3.9, 4.2},
  {0.9, 3.8, 3.9},
  {-0.3, 2.3, 3},
  {-0.7, 1.3, 2.4},
  {-0.8, 0.7, -0.3},
  {-1.3, -0.4, -1.5},
  {-0.9, -0.3, -2.1},
  {-0.9, -0.6, -2.3},
  {-1.3, -0.6, -2.3},
  {-1.7, -0.3, -2},
  {-1.8, -0.4, -2.1},
  {-1.9, -0.5, -2.4},
  {-2, -0.4, -2.1},
  {-2.3, -0.6, -1.9},
  {-2.6, -0.7, -1.6},
  {-2.3, -1, -1.7},
  {-2.4, -1.2, -1.6},
  {-2, -1.2, -1},
  {-1.6, -0.5, 0.2},
  {-0.7, 0.9, 1.2},
  {1, 2.2, 3.9},
  {2.8, 4.4, 5.7},
  {4.2, 5.6, 7},
  {4.6, 7, 7.4},
  {5, 7.6, 7.2},
  {4.2, 7.2, 7.1},
  {2.9, 5.7, 6},
  {1.3, 4.2, 4.5},
  {0.5, 2.6, 2.7},
  {-0.4, 2.6, 1.5},
  {-0.5, 2, 0.3},
  {-0.6, 1.6, 0},
  {-0.2, 1.4, -0.7},
  {-0.2, 0.9, -0.6},
  {-0.3, 0.8, -1.1},
  {0, 0.9, -0.7},
  {0.2, 1.2, -0.7},
  {0.5, 1.3, -0.2},
  {0.1, 1.5, 0},
  {0.2, 1, 0},
  {0, 0, 0.2},
  {-0.3, 0.3, 0.3},
  {0, 0.6, 0.6},
  {1.8, 2.9, 1.2},
  {2.9, 4.7, 3.8},
  {5.4, 6.8, 6.5},
  {6.5, 8.4, 8.3},
  {6.4, 6.2, 9.2},
  {4.8, 6, 6.8},
  {1.4, 5.9, 5.2},
  {1.9, 5.3, 4.8},
  {1.2, 3.9, 3.3},
  {2.3, 3.3, 2.1},
  {2.5, 2.9, 1.4},
  {2.4, 2.6, 1.3},
  {1.3, 2.1, 1.2},
  {0.5, 2.2, 0.4},
  {-0.4, 1.3, -0.3},
  {-0.8, 1.8, -1.5},
  {-0.4, 1, -2},
  {-1.2, 0, -1.8},
  {-1.4, -0.3, -1.8},
  {-1.1, -0.1, -1.6},
  {-1.4, -0.6, -2.5},
  {-1.4, -0.3, -2.8},
  {-0.5, 0.2, -2.5},
  {1.7, 1.8, 0.1},
  {2.8, 4.4, 3.2},
  {5.1, 6.6, 6.3},
  {5.6, 7.4, 8.6},
  {6.3, 8.3, 9.2},
  {5.5, 8.8, 8.4},
  {4.8, 8.4, 7.4},
  {3.8, 7.6, 7.3},
  {3, 7.8, 6.9},
  {2, 6.2, 4.5},
  {0.1, 4.1, 2.3},
  {-0.1, 3.1, 0.9},
  {-0.6, 2.1, -0.7},
  {-0.6, 1.3, -1.5},
  {-0.8, 1.2, -2},
  {-1.5, 0.6, -2.6},
  {-1.8, -0.1, -3},
  {-1.9, -0.9, -3.5},
  {-2.2, -0.7, -4},
  {-1.3, 0.1, -4},
  {-0.5, 0, -3.1},
  {-0.8, 0.2, -2.2},
  {-1.4, -0.3, 2.7},
  {-2.2, -1.2, 2.3},
  {-2.2, -1.4, 2},
  {-1.6, -1.3, 2},
  {-1.7, -1.3, 2.3},
  {-2.1, -1.1, 2.3},
  {-2.4, -0.7, 1.9},
  {-2.7, -0.7, 1.9},
  {-2.8, -1.1, 1.6},
  {-3.1, -1.6, 1.3},
  {-3.4, -2.3, 1},
  {-4, -3, 0.4},
  {-4.5, -3.4, 0},
  {-5.3, -3.6, -0.3},
  {-5.5, -3.9, -0.6},
  {-5.4, -4, -0.6},
  {-5.7, -4.2, -0.7},
  {-5.4, -4.5, -0.6},
  {-5.9, -4.6, -1},
  {-6.4, -4.7, -1.2},
  {-7.5, -4.7, -2},
  {-7.8, -4.7, -3.4},
  {-7.5, -4.6, -4.6},
  {-6.4, -4.4, -4.1},
  {-5.5, -4.1, -4.2},
  {-3.7, -3.3, -2.9},
  {-2, -3, -1.2},
  {-0.1, -1.1, 1},
  {1.6, 0.8, 3.1},
  {3.3, 2.5, 5.4},
  {4.5, 4.2, 7.4},
  {5.8, 5.6, 8.8},
  {6.2, 6.5, 10.3},
  {6.2, 6.8, 10.5},
  {3.9, 5.9, 6.6},
  {1.2, 3.7, 3.3},
  {0.2, 3.2, 1.7},
  {-0.1, 2.3, -0.2},
  {-0.8, 1.9, -1.3},
  {-1.1, 1.2, -2},
  {-1.9, 0.6, -2.6},
  {-1.8, 0.1, -3.3},
  {-2.5, -0.5, -3.8},
  {-3.4, -0.5, -4.3},
  {-4.3, -1.3, -4.7},
  {-4.3, -1.4, -5.1},
  {-4.1, -1.8, -5.2},
  {-4.3, -1.7, -5.8},
  {-4.1, -1.4, -5.5},
  {-0.8, -0.7, -4.9},
  {1.9, 1.7, -1.5},
  {2.8, 4.4, 1.9},
  {3.5, 6.2, 5.4},
  {4.8, 8.4, 7.2},
  {5.5, 9.4, 7.2},
  {4.8, 9.8, 7.8},
  {4.6, 9.5, 7.8},
  {3.8, 7.4, 7.1},
  {2.2, 5.8, 6.1},
  {0.6, 4.1, 4.5},
  {0.3, 2.9, 1.8},
  {-1.3, 1.8, 0.4},
  {-1.1, 1.1, -0.4},
  {-1.7, 0.6, -1.3},
  {-2.3, 0.4, -1.8},
  {-2.7, 0, -2.4},
  {-3.2, -0.3, -2.7},
  {-3.3, -0.7, -3.2},
  {-3.4, -1.2, -3.5},
  {-3.2, -1.4, -3.7},
  {-2.9, -1.6, -4.1},
  {-2.9, -1.5, -4.3},
  {-2.5, -1.2, -4.3},
  {-0.1, -0.3, -3.4},
  {1.6, 1.5, -0.8},
  {2, 2.7, 2.1},
  {3.5, 4.6, 5},
  {4.8, 6.3, 7.2},
  {5.4, 8, 7.6},
  {5.5, 8.1, 7.1},
  {4.8, 7.4, 6.6},
  {3.2, 6.3, 6.2},
  {2.1, 5.1, 5.7},
  {1.5, 3.7, 5},
  {1.3, 2.9, 2.6},
  {1.2, 2.5, 1.6},
  {0.9, 2.7, 1.4},
  {0.9, 2.8, 1.5},
  {0.7, 2.8, 1.5},
  {0.1, 2.7, 1.6},
  {-0.1, 2.3, 1.8},
  {0.3, 2, 1.7},
  {0.1, 1.8, 1.6},
  {-0.2, 1.7, 1.6},
  {-0.3, 1.7, 1.4},
  {-0.3, 1.7, 1.3},
  {-0.3, 1.8, 1.4},
  {0, 1.7, 1.5},
  {0.7, 1.8, 1.6},
  {0.9, 2.2, 2.4},
  {1.6, 3.2, 3.4},
  {2.3, 4.8, 4.1},
  {2.7, 6.2, 4.9},
  {2.9, 6.2, 5.3},
  {3, 5.8, 5.7},
  {2.3, 5, 5.6},
  {1.2, 4, 4.9},
  {0.2, 2.9, 4.1},
  {-1.3, 1.8, 3},
  {-1.5, 1.6, 1.8},
  {-0.4, 1, 1.6},
  {0, 1.5, 1.8},
  {0.1, 2.1, 1.7},
  {0, 1.8, 1.6},
  {-0.9, 1.8, 1.5},
  {-2.2, 0.5, 1.1},
  {-1.6, 0.2, 0.3},
  {-1.1, 0, -0.5},
  {-1.5, 0.5, -0.8},
  {-1.9, 0.2, -1.3},
  {-0.5, 0.5, -1.1},
  {0.4, 1.4, 0},
  {1.4, 2.8, 1.6},
  {2.8, 4.3, 4.5},
  {4.1, 5.5, 7},
  {5.7, 7.1, 8.9},
  {6, 8.5, 9.5},
  {6, 9.3, 9.2},
  {4.9, 8.4, 8.1},
  {3.8, 7, 7.4},
  {2.4, 5.4, 6.5},
  {1.5, 4, 5.6},
  {-0.3, 3.3, 3.4},
  {-0.3, 2.4, 2.1},
  {-0.1, 2.3, 2},
  {0.4, 3, 2.3},
  {0.8, 3.2, 2.5},
  {-0.9, 2.9, 2.6},
  {-0.1, 2.7, 2.7},
  {0.3, 2.6, 2.6},
  {0.1, 2.3, 2.8},
  {-0.4, 2.1, 3},
  {-0.2, 1.7, 2.8},
  {0, 1.7, 2.5},
  {0, 1.8, 2.5},
  {0.2, 2.2, 2.5},
  {0.1, 2.3, 3},
  {0.3, 2.7, 3.4},
  {0.8, 3.7, 3.7},
  {1.4, 4.4, 4},
  {2.3, 5, 4.7},
  {3.3, 5.7, 5.4},
  {3, 5.9, 6.2},
  {3.1, 5.5, 6.5},
  {2.2, 4.4, 6.4},
  {0.3, 3.5, 5.1},
  {0.1, 2.5, 3.7},
  {-0.7, 1.7, 3},
  {-0.4, 0.7, 1.9},
  {0.6, 0.7, 0.6},
  {-0.2, 0.9, 0.4},
  {-1, 1.7, 0.6},
  {-0.8, 1.5, 0.7},
  {-0.4, 1.4, 0.6},
  {-0.3, 1.4, 0.7},
  {-0.4, 1.3, 0.8},
  {-0.1, 1.1, 0.8},
  {-0.2, 1.1, 0.7},
  {0.2, 1.4, 0.9},
  {1, 1.7, 1.9},
  {1.3, 3.8, 3.5},
  {2.3, 5.4, 5.4},
  {4.5, 6.3, 7.7},
  {5.4, 7.4, 9.1},
  {6.2, 8.7, 10.3},
  {6.5, 9.8, 10.9},
  {6.8, 9.9, 10.1},
  {6.8, 9.4, 8.9},
  {3.7, 8.1, 8},
  {1.3, 5.7, 6.5},
  {-0.2, 4, 4.7},
  {-0.6, 3.3, 2.8},
  {-0.8, 2.5, 1},
  {-1.3, 1.9, 0},
  {-1.3, 1.4, -0.6},
  {-1.6, 1, -1.2},
  {-1.6, 1.3, -1.5},
  {-2.1, 0.7, -1.8},
  {-1.9, -0.1, -2},
  {-1.8, -0.3, -2.3},
  {-2.3, -0.5, -2.7},
  {-1.6, -0.3, -2.8},
  {-1, 0.2, -2.6},
  {1.6, 0.7, -1.5},
  {3.5, 2.5, 1},
  {4.5, 4.4, 4.3},
  {5.8, 6.7, 7.6},
  {6.8, 8.4, 9.7},
  {7.4, 10, 10.1},
  {7.8, 10, 9.2},
  {6.9, 9.1, 8.9},
  {6.1, 7.9, 9},
  {4.6, 6.9, 8.7},
  {3.5, 6, 7.5},
  {3.1, 5.2, 5.3},
  {2.9, 4.2, 3.7},
  {2.6, 3.6, 2.6},
  {2.5, 4.1, 1.8},
  {2.2, 4.2, 1.9},
  {0.8, 4.5, 1.6},
  {-0.2, 3.8, 1.9},
  {-0.4, 3.2, 2.2},
  {-0.9, 2.9, 2.2},
  {-0.9, 3.1, 2.3},
  {-0.3, 2.8, 2.3},
  {0.5, 2.7, 1.9},
  {1.6, 2.6, 1.8},
  {2.7, 4, 3},
  {3.5, 4.4, 4.6},
  {3.5, 4.4, 6.2},
  {3.6, 5.5, 7.9},
  {3.5, 6.4, 9.2},
  {3.3, 6.8, 8.6},
  {3.2, 6, 6.6},
  {2.9, 5.2, 6.1},
  {2.6, 4.5, 5.9},
  {2.4, 3.8, 5.4},
  {2.4, 3.3, 4.9},
  {2.2, 3.3, 4.5},
  {2.3, 3.3, 4.3},
  {2.2, 3.3, 4},
  {2.2, 3.2, 3.9},
  {2.4, 3.1, 3.8},
  {2.3, 3.1, 3.7},
  {2, 3.1, 3.5},
  {1.9, 3, 3.3},
  {1.3, 2.9, 3.1},
  {1, 3.1, 2.8},
  {0.9, 3.3, 2.7},
  {0.9, 3.7, 2.4},
  {2, 4.4, 2.7},
  {3.7, 4.6, 3.1},
  {5.1, 6.4, 3.3},
  {7.2, 7.7, 4.3},
  {8.7, 9, 7.9},
  {10, 11.2, 12.2},
  {9.8, 12.3, 14.2},
  {10.2, 13, 14.6},
  {10.1, 13.5, 14.4},
  {10, 13.4, 12.5},
  {8, 12.5, 11.2},
  {5.5, 10.1, 9.8},
  {4, 8.2, 7.6},
  {3.9, 7.4, 5.9},
  {3.7, 7.1, 4.4},
  {4.2, 6.4, 3.7},
  {5, 6, 3.5},
  {4.8, 5.6, 3.4},
  {4.4, 4.7, 2.7},
  {4.4, 4.7, 2.1},
  {3.7, 4.7, 1.4},
  {3.2, 4.4, 1.1},
  {3.8, 3.9, 0.6},
  {3, 3.3, 0.1},
  {4.8, 3.5, 0.2},
  {5.9, 4.6, 1.3},
  {7.2, 7.2, 4},
  {7.6, 8.7, 7.4},
  {9.1, 10.7, 11.5},
  {9.3, 12.2, 13},
  {8.9, 13, 12.6},
  {9.4, 12.6, 12.4},
  {8.9, 11.2, 12.6},
  {8.3, 10, 11.7},
  {7.3, 9.8, 10.8},
  {6.5, 8.3, 10.3},
  {5.7, 7.6, 9.7},
  {5.7, 7.2, 8.3},
  {4.2, 7.4, 7.7},
  {3.2, 6.4, 6.3},
  {3.8, 5.6, 4.7},
  {5, 6.4, 4.8},
  {5, 6.6, 5.4},
  {5, 6.1, 5.6},
  {5, 5.6, 5.4},
  {4.9, 6.3, 5.2},
  {4, 5.8, 4.8},
  {4.1, 5.5, 4.6},
  {5, 6.1, 4.7},
  {5.5, 6.8, 6.1},
  {5.4, 7.6, 7.3},
  {5.4, 8, 8.1},
  {4.1, 7.1, 8.2},
  {2.2, 5.7, 7},
  {2.5, 4.9, 6.4},
  {3.3, 5.2, 6.4},
  {3.4, 5.3, 6.3},
  {3.6, 5.1, 6.5},
  {3.7, 5, 6.8},
  {3.3, 5.1, 6.5},
  {3, 5.1, 6.1},
  {2.6, 4.8, 5.8},
  {2.2, 4.7, 5.7},
  {2.3, 4.6, 5.4},
  {2.5, 4.5, 5.3},
  {2.7, 4.5, 5.1},
  {2.5, 4.2, 5.2},
  {2.8, 4.2, 4.9},
  {2.4, 4, 4.7},
  {2.3, 3.7, 4.4},
  {1.6, 3.7, 4},
  {1.1, 3.4, 3.8},
  {2.3, 4.3, 3.9},
  {4.9, 5.2, 4.9},
  {6.2, 6.1, 6.3},
  {7.4, 7.4, 8},
  {8.5, 9.1, 10.6},
  {9.3, 10.9, 13.2},
  {10.1, 12.3, 13.5},
  {9.9, 13.4, 13.4},
  {9.3, 13, 13.3},
  {8.2, 11.3, 12.5},
  {6.9, 10.5, 11.8},
  {6.1, 9.1, 11.1},
  {5.9, 8.1, 10.1},
  {5.8, 7.4, 8.3},
  {5.8, 7, 7.3},
  {5.8, 6.4, 6.9},
  {5.8, 6.2, 7},
  {5.9, 6.4, 7.1},
  {5.9, 6.3, 7},
  {5.7, 6.7, 6.9},
  {5.6, 6.3, 6.8},
  {5.4, 5.9, 6.7},
  {4.9, 6.1, 6.4},
  {4.3, 6.2, 6.3},
  {5.3, 6.8, 6.6},
  {6, 7.3, 7.3},
  {6.8, 7.5, 8.4},
  {8.1, 8.6, 10.1},
  {9.6, 10.1, 12.1},
  {11, 11.9, 14.2},
  {12.4, 13.9, 16.2},
  {12.9, 15.6, 16.9},
  {11.9, 15.3, 15.4},
  {9.9, 13.5, 14.5},
  {8.9, 11.9, 13.5},
  {8.5, 10.7, 12.4},
  {8.3, 10, 10.8},
  {8.3, 9.5, 9.9},
  {8.1, 9.3, 9.6},
  {7.9, 9.4, 9.3},
  {7.5, 9.3, 9.2},
  {7.2, 8.5, 9.2},
  {6.8, 8.6, 9.1},
  {6.8, 8.3, 8.9},
  {6.7, 8.5, 8.7},
  {6.6, 8.2, 8.6},
  {6.4, 7.6, 8.5},
  {6.2, 7.8, 8.4},
  {6.5, 7.9, 8.5},
  {6.5, 7.8, 8.6},
  {6.7, 8, 9},
  {6.8, 7.8, 9.5},
  {8.1, 7.8, 10.1},
  {8, 8.1, 10.4},
  {8.5, 8.3, 10.8},
  {8.9, 8.7, 11.4},
  {9.4, 9.5, 11.3},
  {9.5, 9.9, 11.4},
  {9.4, 9.4, 11.1},
  {9.1, 9.2, 10.7},
  {8.9, 9.1, 10.2},
  {8.7, 9, 9.5},
  {8.4, 8.9, 8.9},
  {8, 8.7, 8.5},
  {7.6, 8.6, 8.2},
  {7.4, 8.4, 8.2},
  {6.8, 8.2, 8.1},
  {6.7, 8, 8},
  {6.5, 7.8, 8},
  {6.4, 7.6, 7.8},
  {6.7, 7.7, 7.8},
  {7.2, 7.7, 7.8},
  {7, 7.7, 7.9},
  {6.9, 7.6, 8.1},
  {6.5, 7.9, 8.2},
  {6.6, 8.3, 8.7},
  {7.1, 8, 9.1},
  {7.1, 7.8, 9.2},
  {7.4, 7.9, 9.4},
  {7.5, 7.8, 9.3},
  {7.5, 7.8, 9.2},
  {7.2, 7.7, 9.3},
  {7.3, 7.9, 9.2},
  {7.2, 8, 9},
  {6, 7.6, 8.9},
  {5.5, 5.6, 8.6},
  {4.3, 4.9, 7.5},
  {1.3, 4.8, 5.6},
  {1.1, 4.5, 4.7},
  {1.3, 4.2, 4.3},
  {1.7, 4.3, 4.2},
  {1.7, 4.1, 3.7},
  {1.8, 3.7, 3},
  {1.3, 3.2, 2.6},
  {1.2, 2.8, 2},
  {1.2, 2.4, 2.5},
  {2.1, 3.2, 2.9},
  {4.3, 3.8, 3.2},
  {6.9, 5.9, 4.4},
  {8, 8.7, 6.8},
  {8.8, 9.7, 10.1},
  {10, 11, 12},
  {11.2, 12.5, 14},
  {11.8, 13.2, 15.5},
  {11.6, 14, 15.3},
  {11.2, 14.1, 15},
  {9.4, 13.2, 13.7},
  {8.2, 9.5, 11},
  {5.4, 7.9, 8},
  {4.8, 7.3, 6},
  {5.1, 7, 4.7},
  {5, 6.2, 3.6},
  {4.4, 5.5, 2.6},
  {3.2, 4.7, 1.7},
  {3.3, 3.9, 1.2},
  {1.7, 3.6, 0.4},
  {1.6, 3.3, 0.1},
  {2, 3, -0.2},
  {2.6, 2.9, -0.3},
  {2.2, 3, -0.2},
  {3.7, 4.3, 0.4},
  {5.1, 4.8, 1.9},
  {7, 4.5, 4.1},
  {8.2, 5.7, 6.8},
  {9, 7.3, 9.9},
  {9.6, 9.2, 12.6},
  {10.5, 10.9, 14.7},
  {11, 11.8, 13.9},
  {10.1, 11.9, 13.9},
  {9.4, 11.6, 13},
  {9.2, 11.5, 13.2},
  {7, 10, 11.5},
  {6.6, 9, 9.3},
  {5.6, 8.5, 7.8},
  {5.3, 8.2, 6.6},
  {5.8, 7.8, 6.4},
  {5.5, 7.2, 6.1},
  {4.5, 6.5, 5.9},
  {4.1, 6.2, 5.2},
  {4.3, 5.9, 4.3},
  {4.5, 6.3, 4.3},
  {4.7, 6.6, 4.5},
  {5.4, 6.3, 5},
  {5.4, 6.1, 5.3},
  {6.2, 6.3, 5.7},
  {7.2, 7.1, 6.8},
  {8.8, 8.3, 8.8},
  {9.6, 10.8, 11.5},
  {11.4, 12.5, 14.1},
  {12.1, 13.8, 16},
  {13.3, 15.2, 16.6},
  {13.8, 16, 16.8},
  {12.4, 16.2, 16.9},
  {13, 14.9, 17.2},
  {12.3, 14.6, 17.2},
  {11.2, 13.2, 15},
  {8.7, 11.6, 12.4},
  {8, 10.6, 10.4},
  {9.6, 9.8, 8.8},
  {9.5, 9.7, 7.7},
  {9.2, 9.9, 7},
  {8.9, 9.7, 7},
  {8.6, 8.7, 7.2},
  {8, 8.6, 6.7},
  {7.6, 8.2, 7.1},
  {7.3, 8.1, 7},
  {7.2, 7.8, 6.8},
  {7.3, 6.7, 6.4},
  {7.4, 8.1, 6.8},
  {7.6, 8.6, 7.6},
  {8, 9.9, 9},
  {9.8, 11.2, 11.1},
  {10.2, 12.4, 13.8},
  {10.5, 13, 14.5},
  {10.7, 12.5, 13.5},
  {10.4, 12.2, 14.2},
  {10.5, 12.1, 14.5},
  {10.5, 11.9, 14},
  {9.7, 11.5, 13.5},
  {8.4, 10.9, 12.5},
  {8.2, 10.3, 11.8},
  {7.9, 9.9, 11.5},
  {6.2, 9.2, 10.9},
  {5.5, 8.1, 9.9},
  {4.9, 7.7, 8.9},
  {4.8, 7.5, 8.4},
  {5, 7, 8},
  {4.6, 7, 6.8},
  {4.6, 6.7, 5.8},
  {4.8, 7.2, 5.1},
  {4.4, 7.2, 4.7},
  {5.3, 7, 4.1},
  {6.2, 7.2, 4.4},
  {9.3, 8.6, 6.4},
  {10.7, 10.1, 9.7},
  {11.9, 13, 13.5},
  {12.9, 14, 16.5},
  {14, 15.6, 18.8},
  {14.9, 17.2, 18.9},
  {14.3, 17.4, 18.8},
  {13.6, 16.4, 17.5},
  {11.5, 15.2, 15.8},
  {10, 13.6, 14.5},
  {9.7, 12.2, 13.8},
  {9.2, 11, 12.1},
  {9, 10.1, 10.1},
  {7, 9.2, 8.5},
  {6.4, 8.5, 7.4},
  {6.4, 8.3, 6.6},
  {6.3, 7.8, 6.1},
  {6.4, 7.4, 5.5},
  {6.2, 6.9, 5},
  {5.9, 6.9, 4.9},
  {5.6, 6.5, 4.6},
  {5.4, 6.6, 4.4},
  {5.5, 6.8, 4.6},
  {7.6, 7.6, 5.5},
  {8.1, 8, 6.8},
  {9.1, 8.7, 8.4},
  {9.4, 9.6, 10.3},
  {11, 8.8, 12.7},
  {11.8, 6.3, 14.1},
  {9.5, 8.6, 12.2},
  {5.5, 10.9, 10.2},
  {7.2, 12.2, 12.3},
  {8.6, 12.1, 13.3},
  {7.3, 11.9, 12.7},
  {7.5, 9.8, 10.6},
  {6.4, 8.4, 8},
  {6.7, 8.2, 6.3},
  {5.7, 7.3, 5},
  {4.5, 6.5, 3.7},
  {2.8, 6, 2.7},
  {2.2, 5.3, 1.9},
  {2, 4.7, 1.2},
  {1.7, 3.9, 0.5},
  {1.3, 3.7, 0.1},
  {0.7, 3, -0.4},
  {0.3, 2.6, -0.8},
  {0.5, 2.8, -0.9},
  {2.7, 3.2, -0.7},
  {6.9, 5, 1.4},
  {7.8, 7.1, 5.8},
  {9.5, 9.3, 9.7},
  {10.1, 11.4, 13},
  {10.9, 12.7, 14.2},
  {11.2, 13.5, 14.4},
  {10.8, 13.8, 14.1},
  {10.7, 13.4, 14.4},
  {10.2, 12.8, 14.1},
  {9.4, 11.9, 13.3},
  {8.3, 10.3, 12.3},
  {6.5, 8.8, 10.8},
  {5.2, 8.9, 8},
  {6.7, 8.1, 6.2},
  {6.3, 7.9, 5.1},
  {6.5, 7.8, 4.8},
  {5.7, 7.5, 5.1},
  {5.7, 7.3, 5.4},
  {5.1, 5.8, 5},
  {5, 5.6, 4.9},
  {4.8, 5.7, 4.8},
  {5.4, 5.4, 4.7},
  {5.6, 5.6, 4.8},
  {5.8, 6.4, 5},
  {6.2, 6.8, 5.6},
  {6.1, 6.2, 6.3},
  {6.3, 6.8, 7.1},
  {4.9, 7.2, 8},
  {2.4, 5.6, 7.8},
  {3, 3.9, 6.2},
  {2.8, 3.7, 6},
  {2.9, 3.6, 5.7},
  {2.9, 3.6, 5.4},
  {3.1, 3.6, 5.2},
  {3.7, 3.7, 5.2},
  {3.7, 3.7, 5.1},
  {3.6, 3.7, 5.1},
  {3.8, 3.7, 4.9},
  {3.7, 3.8, 4.8},
  {3.6, 3.9, 4.8},
  {3.6, 3.8, 4.8},
  {3.4, 3.8, 4.7},
  {3.1, 3.9, 4.8},
  {2.8, 3.9, 4.7},
  {2.6, 4, 4.7},
  {2.5, 3.6, 4.8},
  {2.1, 3.5, 4.7},
  {2, 3.6, 5},
  {1.8, 4, 5.3},
  {1.7, 4.7, 5.7},
  {2.2, 5.6, 7.2},
  {2.3, 6.2, 8.6},
  {3.1, 6.5, 9},
  {4.1, 7.2, 8.9},
  {3.6, 8.4, 10.6},
  {3.7, 7.6, 10.4},
  {4.3, 7.3, 9.1},
  {4.6, 6.7, 8.6},
  {3.3, 5.2, 7.9},
  {2.1, 3.2, 6},
  {1.7, 2.4, 5.7},
  {1.6, 1.9, 5.6},
  {1, 1.2, 5.4},
  {0.5, 0.8, 4.8},
  {0, 0.9, 3.9},
  {0.3, 0.8, 4.1},
  {0.1, 0, 4.2},
  {0.4, -0.4, 4.1},
  {0.6, -0.3, 3.8},
  {0.7, -0.3, 3.5},
  {0.4, -0.4, 3.6},
  {0, 0.2, 3.9},
  {-0.1, 1.5, 4},
  {0.4, 4, 4.5},
  {1.5, 5.3, 6.4},
  {3.5, 6.9, 8.5},
  {4.6, 8.6, 9.8},
  {6.4, 9.7, 11.1},
  {7.1, 10.4, 11.9},
  {7.5, 10.5, 10.8},
  {7.6, 10.5, 10.7},
  {5.4, 9.6, 9.7},
  {3.5, 7.7, 8.3},
  {1.9, 5.7, 6.9},
  {1.2, 5.1, 5.1},
  {0.8, 4.1, 3.7},
  {0.6, 3.5, 2.6},
  {0.4, 3.1, 1.8},
  {0.4, 2.3, 1},
  {-0.3, 1.9, 0.4},
  {-0.4, 1.4, 0},
  {-0.6, 1.3, -0.4},
  {-0.6, 1, -0.7},
  {-0.6, 1.1, -1},
  {-0.6, 1.3, -1},
  {2.4, 1.9, -0.8},
  {5.1, 3.4, 1.5},
  {6.1, 5.4, 5.4},
  {7.2, 7.8, 9.4},
  {8.7, 10, 12.2},
  {10, 11.8, 14.5},
  {10.7, 13.3, 14.6},
  {11.2, 14, 14.3},
  {11.1, 13.2, 13.2},
  {9.6, 12.4, 12.7},
  {8, 11, 12.3},
  {6.5, 9.3, 10.9},
  {5.9, 8.4, 8.9},
  {5.2, 7.7, 6.7},
  {4.2, 6.8, 5.3},
  {2.9, 7, 4},
  {3.7, 6.3, 3.1},
  {3.2, 4.9, 2.4},
  {2.2, 4.7, 2},
  {2.8, 4.1, 1.5},
  {2.6, 4, 1.5},
  {2.8, 3.9, 1.4},
  {2.3, 3.4, 1.1},
  {3, 4, 1.3},
  {5.4, 5.6, 2.4},
  {6.7, 6, 4.6},
  {8, 7.9, 7.1},
  {8.4, 9.6, 9.4},
  {9.7, 11.1, 11.9},
  {10.2, 11.7, 13.2},
  {10.5, 11.9, 12.9},
  {7.9, 11.7, 12.1},
  {7.9, 11.2, 11.7},
  {8.1, 11, 12},
  {7.6, 9.9, 11.5},
  {7.3, 9.1, 11},
  {7.1, 8.2, 10.2},
  {7.2, 8, 9.3},
  {6.8, 8.2, 8.4},
  {6.5, 8.4, 8},
  {6.4, 8, 7.7},
  {6.4, 7.7, 7.7},
  {6.4, 7.7, 7.5},
  {6.6, 8.2, 7.5},
  {6.5, 8.3, 7.4},
  {6.4, 7.9, 7.3},
  {5.6, 8.1, 7.1},
  {6.7, 8.3, 7},
  {7.5, 8.7, 7.3},
  {7.5, 8.9, 8.1},
  {7.9, 8.9, 8.9},
  {8.1, 8.8, 9.4},
  {7.8, 9, 10},
  {8.8, 9.5, 10},
  {9.2, 10, 10.3},
  {8.3, 10, 10.5},
  {7.8, 9.7, 10.3},
  {7.1, 8.6, 10.1},
  {6.8, 7.7, 9.2},
  {6.2, 7.3, 8.8},
  {6, 7.1, 7.9},
  {6.2, 7, 7.4},
  {6, 6.8, 7.2},
  {5.9, 6, 7},
  {5.6, 5.6, 6.6},
  {5.2, 5.1, 6.3},
  {4.8, 3.8, 5.9},
  {4.1, 3.3, 5.7},
  {3.1, 2.6, 5.5},
  {2, 2.7, 5.4},
  {1.3, 2.5, 5.3},
  {1.4, 1.9, 5.1},
  {2.2, 1.2, 4.5},
  {1.7, 1.3, 4.3},
  {2, 2.1, 4.6},
  {2.2, 3.7, 5},
  {2.8, 5, 6.5},
  {3.4, 6.4, 7.7},
  {4.4, 7.4, 8.4},
  {4.9, 8.2, 9.3},
  {5.6, 8.6, 10.1},
  {5.9, 8.3, 11.2},
  {5.5, 7.1, 10.7},
  {5.2, 6.1, 10.1},
  {5.2, 5.6, 9.4},
  {4.8, 5.2, 8.4},
  {4.3, 4.6, 6.8},
  {2.7, 3.8, 5.1},
  {0.4, 3.4, 3.2},
  {0.2, 3.1, 1.8},
  {-1, 2.4, 1.2},
  {-1, 2.6, 0.6},
  {-1.8, 1.8, 0},
  {-1.2, 1.1, -0.5},
  {-0.5, 1.8, -0.6},
  {0.2, 1.8, -0.3},
  {0.9, 2.5, 0.6},
  {2.1, 2.9, 1.9},
  {2.3, 4.1, 2.9},
  {3.2, 4.1, 4.1},
  {3.4, 5.8, 5.9},
  {5.2, 7, 7.9},
  {6.4, 8.5, 9.8},
  {7.2, 9.5, 10.9},
  {8.2, 10.6, 12},
  {8.8, 11, 12.5},
  {7.6, 10.3, 12.8},
  {6.4, 8.1, 10.8},
  {5, 7.2, 9.7},
  {3.4, 6.8, 8.3},
  {3.2, 5.9, 6.1},
  {2.1, 4.9, 4.3},
  {1.8, 4.2, 2.9},
  {1, 3.4, 1.8},
  {0.4, 2.9, 1},
  {0.3, 2.3, 0.4},
  {0, 2.2, -0.1},
  {0, 1.8, -0.5},
  {-0.1, 1.8, -1},
  {0.9, 1.9, -1.1},
  {4, 3, -0.6},
  {6.1, 5.6, 2.4},
  {7.1, 8.4, 6.1},
  {8.5, 10.3, 10},
  {9.5, 11.4, 12.7},
  {10.5, 11.9, 13.9},
  {11.1, 12.9, 15.3},
  {10.7, 13.9, 15},
  {10.5, 14.1, 14.5},
  {10.3, 14.3, 14.2},
  {9.1, 13, 14.3},
  {8.3, 11.2, 12.5},
  {7.9, 10.1, 9.7},
  {7.5, 8.5, 7.4},
  {5.2, 6.8, 5.9},
  {4.5, 6.3, 4.6},
  {4.2, 5.9, 3.5},
  {3.5, 5.9, 3},
  {3.5, 5.3, 2.5},
  {3.3, 4.7, 1.9},
  {2.9, 4.4, 1.4},
  {2.6, 4.3, 1},
  {2.8, 4, 0.6},
  {3.6, 4.3, 0.7},
  {7.3, 5.1, 1.4},
  {9.2, 7.3, 5.5},
  {10.5, 9.8, 9.6},
  {11.4, 11.5, 13.2},
  {12.9, 13.6, 15.7},
  {14.2, 15.6, 16.5},
  {15.2, 16.6, 16.6},
  {15.1, 16.5, 17.6},
  {15.2, 16.4, 18},
  {13.9, 16.4, 18},
  {13, 15.5, 17.4},
  {12.3, 14.1, 15.8},
  {11.5, 12.5, 13},
  {11.5, 12.3, 10.9},
  {10.6, 12.2, 8.9},
  {10.6, 10.8, 7.8},
  {9.7, 9.5, 6.9},
  {8, 9.1, 6.1},
  {6.7, 8.4, 5.4},
  {6.4, 7.7, 5},
  {5.6, 7.1, 4.4},
  {5.1, 6.6, 4},
  {4.9, 6.6, 3.5},
  {5.8, 7.1, 3.8},
  {7.5, 8.1, 4.8},
  {8.6, 9.4, 7.5},
  {9.3, 10.6, 9.8},
  {11.1, 11.6, 12.8},
  {12, 13, 15.1},
  {11.4, 13, 14.5},
  {10.6, 12.2, 13.1},
  {9.4, 11.1, 13},
  {8.2, 10, 12},
  {7.6, 9, 10.6},
  {7.7, 8.9, 10.2},
  {8, 8.6, 10.1},
  {7.8, 8.3, 9.8},
  {8.5, 8.8, 9.4},
  {8.7, 9, 9.1},
  {8.4, 8.9, 8.9},
  {8, 8.6, 8.8},
  {7.7, 8.4, 8.7},
  {7.4, 8.2, 8.2},
  {7.1, 8.3, 8},
  {7, 8.2, 8.1},
  {7.2, 8.1, 8},
  {7.1, 8.2, 8},
  {7, 8.3, 8},
  {7, 8.5, 8.2},
  {7, 9.2, 8.8},
  {7.4, 9, 9.1},
  {8.3, 10.3, 10.1},
  {9.5, 11.2, 12.1},
  {10.2, 12.4, 13.8},
  {10.8, 13.4, 14.7},
  {11.8, 14.9, 16.4},
  {12.2, 15.4, 16.7},
  {12.4, 14.8, 16.3},
  {11.1, 14, 15.6},
  {9.6, 13.2, 14.8},
  {8.7, 11.2, 13.2},
  {8.9, 9.9, 11.5},
  {9.1, 9.8, 10.9},
  {8.9, 10.2, 10.3},
  {9.2, 10.2, 9.4},
  {9.3, 9.8, 9.4},
  {7.6, 9.5, 9.5},
  {7.2, 9.2, 9},
  {7.8, 8.4, 8.8},
  {7, 8.2, 7.9},
  {6.9, 8.3, 6.7},
  {7.8, 8.4, 6.5},
  {8.2, 8.4, 7.5},
  {9, 10.1, 9.6},
  {10.5, 10.4, 11.6},
  {11.5, 12.1, 13.7},
  {11.6, 13.8, 16.5},
  {11.6, 15.6, 16},
  {12.3, 15.7, 16},
  {12.7, 15.7, 16.4},
  {12.2, 15.2, 16.6},
  {11, 14.8, 16.6},
  {10.7, 14.4, 15.5},
  {10.3, 13.2, 14.7},
  {9.4, 11.3, 13.6},
  {8.3, 10.9, 11.8},
  {7.6, 10.1, 9.9},
  {7.3, 9.8, 8.6},
  {7.8, 8.7, 7.4},
  {8, 9.2, 6.9},
  {7.8, 9.7, 7.2},
  {7.8, 9, 7.5},
  {7.3, 8.7, 7.5},
  {7, 8.5, 7.6},
  {6.8, 8.6, 7.4},
  {7, 9, 7.4},
  {7, 9.2, 7.9},
  {6.9, 9.6, 8.5},
  {7.4, 9.9, 9.1},
  {8.4, 10.8, 9.7},
  {10.4, 12.2, 11.3},
  {12.4, 13.7, 14.2},
  {12.8, 14.1, 16.7},
  {11.9, 13.9, 17.9},
  {11.1, 13.1, 17.3},
  {11.4, 13, 16.2},
  {10.6, 13.4, 16.1},
  {10, 11.9, 15.5},
  {9.4, 10.1, 14.5},
  {8.3, 9.9, 12.9},
  {7.1, 9.3, 10.6},
  {7.3, 8.7, 9.2},
  {7.1, 8.3, 7.9},
  {6.6, 8.1, 6.7},
  {6.1, 8.6, 6},
  {6.7, 8.3, 5.3},
  {6.5, 8, 4.8},
  {5.7, 7.7, 4.6},
  {4.8, 7.6, 4.2},
  {6, 8.5, 3.7},
  {7.8, 9.7, 4.3},
  {8.7, 10.9, 6.7},
  {10.3, 13.2, 9.1},
  {10.8, 13.1, 13.5},
  {11.8, 14.3, 15.9},
  {12.7, 14.9, 16.9},
  {13.8, 15.1, 16.8},
  {13.7, 15.4, 17.6},
  {13.1, 16, 17.2},
  {11.4, 15.4, 16.2},
  {9.6, 13.4, 15.6},
  {9.1, 12.2, 14.2},
  {8.9, 11.2, 13},
  {7.6, 10.7, 12},
  {6.8, 10.3, 10.2},
  {7.1, 9.6, 9.4},
  {7.9, 8.7, 9.4},
  {7.7, 8.4, 9.2},
  {7, 8.4, 9.2},
  {5.8, 7.6, 8.4},
  {5.8, 7, 6.9},
  {5.2, 6.3, 5.8},
  {4, 6.1, 4.9},
  {5.3, 6.3, 4.7},
  {8.2, 7.4, 5.8},
  {9.5, 9.3, 9.8},
  {10.6, 11.4, 12.9},
  {12, 13.1, 15.5},
  {13.7, 15.1, 17.9},
  {14.8, 17.5, 19.6},
  {15, 18.2, 18.3},
  {14.8, 17.9, 19.6},
  {14.6, 18.1, 18.6},
  {13.1, 16.6, 17.9},
  {12.6, 15.7, 17.6},
  {11.8, 14.2, 15.7},
  {9.8, 12.9, 14},
  {8.2, 12, 11.7},
  {7.6, 11.3, 10.1},
  {7.3, 10.8, 8.6},
  {7.6, 10.5, 7.9},
  {7.8, 9.9, 6.9},
  {8.3, 8.8, 6.3},
  {7.7, 8, 5.8},
  {6.7, 7.9, 5.3},
  {6.1, 7.6, 4.6},
  {6.1, 7.4, 4.2},
  {7.2, 8.2, 4.2},
  {10.2, 9.1, 5.2},
  {11.6, 10.3, 9.5},
  {13.4, 12.5, 12.6},
  {14, 14.6, 15.9},
  {14.7, 16.2, 18.8},
  {14.6, 17.8, 19.1},
  {15, 18.6, 19.5},
  {14.9, 18.5, 19.8},
  {15.4, 18.4, 20.4},
  {15.5, 17.5, 17},
  {13.2, 16.8, 16.5},
  {12.5, 15.6, 16.2},
  {11.9, 13.6, 13.6},
  {9.8, 12.6, 11.4},
  {9, 11.2, 9.6},
  {8.3, 10, 8.5},
  {7.9, 9.3, 7.6},
  {7.2, 8.7, 6.9},
  {7.1, 8.2, 6.1},
  {7.2, 8.4, 5.4},
  {6.7, 7.9, 4.7},
  {6.3, 7.4, 4.2},
  {6.4, 7.2, 3.8},
  {7.9, 7.6, 3.6},
  {10.7, 8.9, 5.4},
  {11.6, 11.7, 9.5},
  {13.3, 13.1, 13},
  {15, 14.5, 16.9},
  {16.1, 16.8, 19.8},
  {16.9, 19, 21.5},
  {17.2, 20.2, 21.2},
  {15.6, 20.4, 20.7},
  {15.1, 19.3, 19.4},
  {14.1, 18.6, 19.6},
  {14.5, 17.5, 19.7},
  {13.5, 16.6, 18.8},
  {11.1, 14.5, 15.8},
  {9.8, 14.2, 13.1},
  {9.5, 13.8, 11.2},
  {9.5, 12.9, 10.1},
  {8.7, 11.9, 8.9},
  {8.9, 11.4, 7.9},
  {8.2, 10.3, 7.2},
  {7.6, 9.3, 6.5},
  {7.4, 8.7, 5.8},
  {7.4, 9, 5.2},
  {7.2, 9.1, 4.5},
  {9, 9.4, 4.9},
  {12.6, 10.3, 7.3},
  {14.4, 12, 10.9},
  {15.2, 14.1, 14.6},
  {15.8, 16.4, 17.7},
  {16.6, 18.5, 20.4},
  {17.3, 19.5, 21.4},
  {17.2, 20.2, 21},
  {16.3, 20, 21.1},
  {16.2, 19.5, 20.5},
  {16.3, 18.9, 19.7},
  {15.8, 18.6, 20.3},
  {14, 17.1, 18.8},
  {11.2, 15.1, 16.2},
  {11, 14, 13.6},
  {10.7, 13.3, 12},
  {9.5, 13.8, 10.8},
  {9.1, 12.4, 9.8},
  {9.4, 11.1, 8.8},
  {8.8, 10.5, 7.9},
  {8.5, 10, 7.3},
  {8, 9.3, 6.5},
  {7.8, 8.7, 6},
  {7.8, 8.7, 5.5},
  {10.2, 9.1, 5.5},
  {12.5, 10.2, 7.7},
  {13.8, 12.7, 11.7},
  {15.2, 14.4, 15.2},
  {16.4, 16.4, 18.4},
  {17, 18.6, 20.8},
  {17.1, 19.9, 20.8},
  {16.7, 19.8, 20.7},
  {17, 19.7, 21.1},
  {16.8, 20.2, 21},
  {16.3, 19.2, 20.5},
  {16.4, 17.9, 20.6},
  {15.3, 17.1, 19.7},
  {13.1, 15.4, 17.3},
  {11, 15.3, 14.1},
  {10.3, 14.8, 12.1},
  {11.2, 13.8, 11},
  {12, 13, 9.7},
  {11.4, 12.4, 9},
  {9.7, 11.5, 8.2},
  {9.3, 10.6, 7.8},
  {9.9, 10.1, 7.8},
  {10, 10.4, 8.4},
  {9.4, 11, 8.7},
  {11, 11.1, 8.4},
  {13.6, 12.4, 10.6},
  {14.6, 13.3, 13.8},
  {15.3, 14.4, 16.6},
  {16.6, 16.3, 19},
  {16.4, 18.3, 20.5},
  {17, 18.6, 20.8},
  {16.3, 18.8, 21.1},
  {16.2, 19.2, 22.6},
  {17, 20.2, 22.1},
  {15.9, 17.9, 21.1},
  {15.3, 16.6, 20.3},
  {14.6, 16, 19.7},
  {13.3, 15.2, 18.1},
  {12.8, 14.9, 16.1},
  {11.9, 14.7, 14.7},
  {11, 14.2, 14.1},
  {11.1, 13.2, 13.3},
  {11.6, 12.7, 12.9},
  {11.5, 12.5, 12.6},
  {11.7, 12.3, 12.2},
  {10.8, 12.1, 12},
  {10.8, 11.8, 11.7},
  {10.6, 11.8, 11},
  {11.3, 12.1, 10.8},
  {11.6, 12.2, 12.1},
  {12.7, 13.9, 13.9},
  {14.3, 15, 15.4},
  {15.8, 17.2, 17.1},
  {16.2, 17.3, 18.6},
  {15.7, 16.5, 19.4},
  {14.9, 13.4, 19.8},
  {12.2, 12.6, 17.9},
  {11.6, 11.3, 14.5},
  {12.4, 12.1, 13.8},
  {12.1, 12.2, 14.1},
  {11.5, 11.3, 13.4},
  {9.8, 10.4, 13.1},
  {8.8, 10.3, 11.8},
  {7.6, 9.8, 10.4},
  {7.5, 9.8, 9.8},
  {7.3, 10.1, 9},
  {7.6, 9.9, 8.3},
  {7.8, 9.8, 7.7},
  {7.1, 9.7, 7.2},
  {6.5, 9.1, 6.5},
  {6.5, 8.7, 5.8},
  {6.2, 8.9, 5.4},
  {8.1, 9.4, 5.7},
  {10.4, 10.6, 7.3},
  {11.4, 11.3, 9.2},
  {11.9, 12.5, 11.7},
  {12.6, 13.4, 14.5},
  {12.5, 14, 16.2},
  {12.8, 14.2, 17.8},
  {12.1, 14.4, 17.9},
  {11.9, 13.9, 16.6},
  {11.9, 14.2, 16.3},
  {11.7, 13.8, 15.5},
  {10.9, 13.2, 15.3},
  {10.4, 12.5, 14.3},
  {9.8, 11.8, 13.6},
  {9.6, 11, 12.8},
  {9.5, 10.5, 12.4},
  {9.2, 10.4, 12},
  {8.9, 10.2, 11.7},
  {8.7, 10.1, 11.7},
  {8.4, 9.9, 11.5},
  {8.3, 9.7, 11.4},
  {8.4, 9.6, 11.3},
  {8.3, 9.5, 11.1},
  {8.4, 9.5, 10.9},
  {8.5, 9.7, 10.9},
  {9, 10.1, 11.1},
  {9.8, 11.7, 11.4},
  {10.9, 12.8, 12.6},
  {11.6, 13.9, 14.9},
  {12.4, 14.9, 16.6},
  {13.2, 15.1, 19.1},
  {11.7, 15.4, 18.1},
  {10.8, 15.4, 15.1},
  {11.6, 16.1, 14.9},
  {11.9, 15.7, 17.4},
  {11.4, 14, 16.6},
  {10.3, 13.2, 15.1},
  {9.7, 12.2, 13.3},
  {9.1, 12, 12},
  {8.5, 11.3, 11.6},
  {8.5, 10.7, 11.3},
  {8.8, 10.6, 11.1},
  {8.5, 10.1, 10.9},
  {8.2, 9.6, 10.8},
  {8.1, 9.8, 10.6},
  {8, 9.5, 10.3},
  {7.9, 9.2, 10.2},
  {8, 8.9, 10},
  {8.4, 9.4, 10},
  {9.1, 9.8, 10.2},
  {9.6, 10.4, 10.9},
  {10.4, 11.5, 12.2},
  {11.4, 12.6, 13.4},
  {11, 14.2, 14.7},
  {10.9, 14.6, 15.7},
  {11.6, 14.6, 16.6},
  {11.9, 14.7, 16.1},
  {11.2, 14, 14.7},
  {11.4, 13.3, 14.6},
  {10.5, 12.8, 16},
  {10.1, 11.9, 14.2},
  {9.3, 10.8, 13.4},
  {9.1, 7.7, 13},
  {8.1, 5.5, 11.1},
  {7, 3.9, 8.9},
  {4.8, 2.7, 7.5},
  {3.1, 2.8, 6.5},
  {1.8, 2.9, 5.9},
  {1.9, 2.4, 5.6},
  {1.7, 2.7, 5.3},
  {1, 2.3, 4.4},
  {0.6, 1.9, 3.5},
  {1.3, 2, 3},
  {2.6, 2.9, 4.1},
  {4.1, 4.2, 5.8},
  {6, 6.1, 8.8},
  {7.4, 8.1, 10.7},
  {9, 9.7, 12.3},
  {10.1, 11.5, 13.6},
  {10.5, 12.8, 15},
  {10.2, 13.4, 14.4},
  {8.7, 13.6, 12.8},
  {7.9, 12.3, 12.4},
  {6.9, 11.1, 12.1},
  {6.4, 9.5, 11.1},
  {5.9, 8.1, 10.3},
  {5.8, 7.8, 9.8},
  {5.1, 7.5, 9.5},
  {4.8, 7.3, 9.2},
  {5, 7.3, 9},
  {4.4, 6.7, 9},
  {3.2, 5.9, 8.7},
  {2.6, 5.7, 8.6},
  {3, 4.9, 8.4},
  {2.9, 4.7, 8},
  {3.1, 5.2, 7.5},
  {4.6, 6.1, 7.5},
  {6.8, 7.1, 8.5},
  {7.6, 8, 10.4},
  {9, 10.4, 12},
  {10.1, 11.1, 14},
  {10.9, 13, 15.7},
  {11.7, 14.5, 14.8},
  {11.7, 14.9, 13.4},
  {11.6, 14.2, 13.5},
  {12.3, 14.2, 13.7},
  {12, 13.7, 14.6},
  {10.4, 12.5, 14},
  {8.8, 11.4, 13.2},
  {8.7, 10.6, 12.6},
  {8.4, 10.2, 11.6},
  {8.1, 10.1, 10.8},
  {8.2, 10, 10.4},
  {8.1, 10.1, 9.9},
  {7.8, 9.9, 9.2},
  {7, 9.1, 9.1},
  {7.5, 8.7, 8.8},
  {7.4, 9.3, 8.8},
  {7.4, 9.1, 8.7},
  {7.5, 9, 8.5},
  {7.7, 9.8, 8.9},
  {7.8, 10.5, 9.3},
  {7.4, 10.5, 9.8},
  {8, 10.9, 10.8},
  {9, 11.8, 11.6},
  {9, 12.9, 12.9},
  {10.2, 13.9, 14.5},
  {11.1, 14.2, 15.9},
  {12.3, 15.7, 17},
  {11.5, 15.5, 15.1},
  {10.8, 14.7, 15.2},
  {10.3, 14.2, 14.7},
  {9.8, 12.8, 13.9},
  {8.8, 11.3, 12.7},
  {9.3, 10.3, 10.6},
  {9.3, 9.5, 9.5},
  {8.1, 9.8, 9.2},
  {7.6, 9.4, 9.3},
  {6.9, 9, 9.5},
  {6.3, 8.3, 8.8},
  {6.2, 8.1, 7.3},
  {5.9, 8.5, 6.7},
  {5.9, 8.7, 6},
  {6.2, 8.3, 5.6},
  {8.4, 8.4, 5.6},
  {10.4, 9.5, 7.5},
  {10.9, 12.2, 10.8},
  {12.4, 13.6, 14},
  {14, 15.4, 17.1},
  {15.3, 17.1, 19.3},
  {16.1, 18.6, 21.2},
  {16.2, 20.1, 20.7},
  {16.7, 20, 19},
  {16.8, 19.7, 19.3},
  {16.4, 19, 19.1},
  {15.2, 17.4, 18.9},
  {13.5, 16.2, 17.6},
  {11.6, 14.4, 16.2},
  {9.5, 13.8, 14.6},
  {8.8, 12.7, 13.2},
  {8.8, 12.8, 12},
  {9.7, 13.1, 11.7},
  {9.1, 13.3, 11.4},
  {9, 12.8, 10.8},
  {8.7, 12.1, 10.3},
  {9.6, 11, 9.9},
  {9.1, 10.1, 9.2},
  {8, 9.4, 8.2},
  {10.8, 10, 8.1},
  {12.6, 11, 9.3},
  {13.7, 13.9, 12.4},
  {13.1, 15.6, 16.5},
  {13.6, 17.2, 19},
  {14.9, 18.5, 20.2},
  {14.9, 18.5, 19.7},
  {14.7, 18.4, 19.6},
  {14.2, 18.3, 19.1},
  {14, 17.9, 19},
  {14.1, 17.6, 18.1},
  {13.7, 16.2, 17.5},
  {13, 15.3, 16.7},
  {12.3, 14.8, 16.3},
  {11.9, 14.5, 15.9},
  {11.6, 13.4, 15},
  {10, 12.5, 14.8},
  {9.1, 11.7, 14},
  {8.8, 11.2, 12.5},
  {8.3, 9.6, 11.8},
  {8.1, 8.6, 11.4},
  {8, 8.3, 11},
  {7.9, 8, 10.6},
  {7.4, 8.1, 10.4},
  {7.4, 8.7, 10.3},
  {7.8, 8.7, 11},
  {8.9, 9.2, 11.8},
  {9.8, 10.2, 12.7},
  {10.4, 9.9, 13.4},
  {10.3, 10.6, 13.5},
  {10.2, 11.9, 14.2},
  {9.8, 11.2, 14.4},
  {9.9, 11, 14.1},
  {9.7, 10.8, 13.9},
  {9.7, 10.7, 13.7},
  {9.6, 10.3, 13.6},
  {9.3, 9.5, 13.1},
  {8.5, 8.9, 12.5},
  {8.3, 8.6, 11.9},
  {8.1, 8.5, 11.3},
  {8.1, 8.6, 11.1},
  {8, 8.6, 10.6},
  {7.7, 8.8, 10.3},
  {7.1, 8.4, 9.8},
  {7.3, 8, 9.3},
  {7, 8, 9.2},
  {6.7, 8.1, 8.9},
  {7.2, 8.2, 8.7},
  {8.5, 8.9, 9.3},
  {9.5, 9.6, 10.6},
  {11.7, 10.7, 12.4},
  {11.5, 11.9, 13.6},
  {11.4, 12.9, 15},
  {12.5, 14.1, 16.1},
  {13.2, 14.8, 17},
  {14.3, 15.4, 18},
  {13.8, 15.2, 18.7},
  {13.7, 13.9, 18},
  {12.6, 13.8, 17.8},
  {12.3, 12.6, 17.3},
  {11.1, 11.7, 15.6},
  {8.6, 10.4, 13.9},
  {7.7, 9.3, 12.3},
  {7.3, 9, 11.2},
  {7.3, 8.8, 9.6},
  {6.6, 8.3, 8.5},
  {6.9, 7.9, 7.5},
  {6, 7.6, 6.6},
  {5.3, 7.2, 6},
  {4.9, 6.7, 5.3},
  {4.6, 6.3, 4.7},
  {5, 6.2, 4.2},
  {8.4, 6.5, 4.7},
  {9.4, 8, 7},
  {10.4, 10.9, 10.4},
  {12, 12.5, 13.5},
  {13.8, 14.2, 16.6},
  {15.2, 15.9, 19.3},
  {16.2, 17.9, 21.1},
  {16.3, 19.5, 20.5},
  {15.9, 19.4, 19.7},
  {15.3, 18.3, 19},
  {14.5, 17.5, 18.3},
  {13.9, 16.6, 18.2},
  {13, 15.7, 17.4},
  {11.9, 14, 16},
  {10.4, 13.3, 13.4},
  {9.4, 13, 11.3},
  {10.3, 12.7, 10.1},
  {9.5, 12.4, 9.8},
  {9.6, 12.2, 9.6},
  {10.1, 11.9, 9.6},
  {9.3, 11.5, 9.5},
  {9.3, 11.1, 9.3},
  {9.7, 11.4, 9.3},
  {9.6, 11.2, 9.5},
  {9.7, 11.4, 9.9},
  {11, 12, 11},
  {11.7, 12.3, 13.4},
  {11.3, 13.6, 14.9},
  {11.2, 14.4, 16.2},
  {11.8, 15.1, 16.1},
  {11.8, 15.6, 15.6},
  {12, 15.9, 16.4},
  {12.3, 16, 15.9},
  {12.4, 15.4, 16.5},
  {12.6, 15.3, 17.2},
  {11.9, 14.4, 16.7},
  {11.2, 13.7, 15.5},
  {10.5, 13, 14.9},
  {10.7, 12.5, 14.2},
  {10.4, 12.4, 13.3},
  {9.3, 12, 12.4},
  {9.4, 10.5, 11.4},
  {9.3, 10.1, 11},
  {8.4, 9.9, 10.7},
  {8.5, 9.6, 10.4},
  {8.2, 9.4, 10.2},
  {7.5, _, 10.2},
  {6.6, 9, 9.9},
  {6.4, 8.1, 9.3},
  {7, 7.7, 8.9},
  {5.1, 7.7, 9.1},
  {3.5, 7.9, 6.8},
  {3.1, 7.4, 6.6},
  {3.6, 6, 6.9},
  {4.4, 6.5, 7.2},
  {6.1, 6.5, 7.6},
  {6.7, 7.3, 8},
  {6.3, 6.9, 8.2},
  {6, 7, 8.2},
  {5.9, 7.3, 8.1},
  {5.8, 7.2, 8.4},
  {6, 6.9, 8.3},
  {6, 6.7, 8.3},
  {5.7, 6.6, 8.2},
  {5.7, 6.4, 8},
  {5.6, 6.1, 7.8},
  {5.5, 6, 7.5},
  {5, 6.1, 7.7},
  {4.3, 6.1, 7.5},
  {4.2, 6.2, 7.5},
  {4.6, 6.1, 7.5},
  {4.8, 6, 7.2},
  {7.6, 6.5, 7.2},
  {8.9, 7.5, 7.3},
  {9.9, 10.6, 7.8},
  {11.6, 12.2, 9.6},
  {12.6, 13.3, 12.9},
  {13.9, 15.7, 17},
  {15, 17.3, 19.3},
  {15.8, 17.5, 20.3},
  {15, 18.7, 20},
  {14.4, 18, 18.9},
  {13.9, 17.1, 17.8},
  {12.6, 16.2, 16.7},
  {11.6, 14.9, 15.4},
  {9.4, 12.9, 14.1},
  {9.1, 12.4, 13.3},
  {9.8, 10.3, 12.3},
  {9.5, 8.8, 11.6},
  {8.5, 8.4, 11.3},
  {7.7, 8.1, 10.6},
  {7.9, 8, 10.2},
  {7.8, 7.7, 9.8},
  {7.4, 7.6, 9.1},
  {7.5, 7.4, 8.8},
  {7.4, 7, 8.7},
  {8.2, 7.4, 9},
  {9.5, 8, 10.3},
  {11.1, 10.1, 12.4},
  {11.6, 12.5, 14.7},
  {12.2, 14.6, 17},
  {14.2, 16.3, 18.8},
  {16.1, 18, 20.6},
  {15.7, 19.3, 20.4},
  {15.3, 19.9, 19},
  {15.2, 19, 18.9},
  {14.8, 18.5, 18.7},
  {13.5, 17.4, 18.1},
  {12.6, 16, 17.2},
  {12.1, 14.2, 16.3},
  {10.9, 12.9, 14.1},
  {10, 12.2, 12.5},
  {9.3, 11.6, 11.5},
  {8.9, 11.1, 11},
  {8.8, 10.5, 11},
  {9, 10.3, 10.6},
  {9.1, 10.1, 10.7},
  {9.2, 10.1, 10.5},
  {9.5, 9.9, 9.7},
  {9.3, 10.2, 9.5},
  {10.7, 10.9, 10},
  {12.6, 11.3, 11.4},
  {14, 13, 13.7},
  {14.7, 15.4, 16.6},
  {15.6, 16.9, 18.8},
  {16.1, 18.1, 19.5},
  {17, 19, 19.9},
  {17, 19.5, 19.6},
  {16.3, 19.2, 19.8},
  {16.2, 19.2, 19.6},
  {16.2, 18.2, 19.6},
  {15.9, 17.8, 20.1},
  {15.1, 16.9, 18.8},
  {13.9, 14.9, 17.8},
  {13.8, 14.4, 15.1},
  {13.5, 14.3, 13.8},
  {11.5, 14, 12.5},
  {10.6, 13.4, 11},
  {10.2, 12, 9.6},
  {9.4, 11.1, 8.6},
  {9, 10.1, 7.8},
  {8.3, 9.3, 7.5},
  {8.6, 9.1, 7.3},
  {9.6, 10.2, 7.5},
  {11.5, 11.1, 8.4},
  {12.8, 12.4, 10.4},
  {14, 13.3, 11.5},
  {15.2, 15, 12.9},
  {15.8, 17, 17.8},
  {16.2, 18.4, 19.4},
  {16.2, 18, 19.5},
  {15.8, 18.6, 19.2},
  {16.1, 18, 19.2},
  {15.9, 18.8, 19.7},
  {15.9, 17.8, 19.5},
  {15, 17.7, 19},
  {14.3, 16.6, 18.4},
  {12.2, 15, 17.4},
  {11, 13.9, 15.1},
  {10.5, 13.4, 13.2},
  {10.8, 13.8, 12.1},
  {11.1, 13.9, 12.1},
  {11.3, 13.7, 11.9},
  {10.6, 13, 11.7},
  {9.7, 11.5, 11.7},
  {9.1, 10.6, 11.2},
  {8.7, 10.2, 11},
  {8.6, 10.1, 11},
  {8.9, 10.4, 11.1},
  {9.7, 10.8, 11.4},
  {10, 11.8, 12.4},
  {11.4, 13.1, 14.3},
  {13.4, 14.5, 15.5},
  {13.9, 15.7, 17.6},
  {14.7, 16.9, 19.8},
  {15.4, 17.6, 20.7},
  {15.3, 18, 19.6},
  {14.9, 17.6, 18.8},
  {15.4, 20, 19.4},
  {14.6, 19.6, 19.4},
  {11.7, 17.8, 17.3},
  {11, 14.6, 15.5},
  {11.3, 13.5, 13.4},
  {10.6, 12, 12.4},
  {9.4, 10, 11.6},
  {8.8, 10.4, 10.5},
  {8.9, 9.3, 9.6},
  {9.2, 8.9, 9},
  {9.8, 8.6, 8.4},
  {9.5, 8.6, 8.1},
  {8.7, 8.1, 7.6},
  {9.3, 8.3, 7.7},
  {10.1, 8.5, 8.7},
  {10.9, 9.9, 9.9},
  {11.3, 12.6, 11.9},
  {12.4, 13.8, 14.1},
  {13.1, 15.6, 16.9},
  {13.2, 17, 18.9},
  {14.4, 17.4, 18.4},
  {15.1, 17.7, 18.5},
  {16, 18.1, 19.8},
  {15.1, 18.1, 19.5},
  {14.5, 17, 18.9},
  {14.1, 16.6, 18.9},
  {13.5, 16.6, 18.6},
  {13, 15.1, 17.2},
  {12.8, 14.2, 15.5},
  {12.2, 13.6, 13.9},
  {11.3, 13, 12.3},
  {9.7, 12.4, 11.4},
  {9.7, 11.8, 10.4},
  {9.4, 11.1, 9.9},
  {9, 10.8, 9.3},
  {8.9, 10.7, 8.9},
  {9.8, 11.1, 9.1},
  {10.6, 11.5, 9.5},
  {12.2, 12, 10.1},
  {14.2, 12.9, 12.3},
  {14.8, 14.9, 14.8},
  {15.6, 15.6, 17.7},
  {16.7, 17.3, 19.9},
  {17.9, 19.8, 22},
  {17.8, 20.3, 21.1},
  {18.1, 20.4, 21.6},
  {17.6, 20.2, 21.2},
  {18.8, 19.8, 21.5},
  {18.8, 20.5, 22.2},
  {17.6, 19.5, 21.6},
  {16.9, 18.8, 21},
  {15.5, 17.5, 20.1},
  {15.6, 16.7, 18.2},
  {15.9, 16.6, 16.9},
  {15.7, 16.5, 15.7},
  {14.4, 15.8, 14.5},
  {12.7, 14.6, 13.5},
  {11.2, 13.6, 12.4},
  {11, 12.9, 11.7},
  {10.8, 12.7, 11.1},
  {10.9, 12.2, 10.6},
  {11.9, 13.1, 10.2},
  {14.5, 14.1, 11.5},
  {14.9, 15.1, 13.7},
  {16.1, 17, 16.4},
  {17.4, 18.4, 19.3},
  {18.9, 20.2, 22.1},
  {19.8, 22.2, 24.4},
  {20.5, 24.3, 25.7},
  {20.9, 24.7, 25.3},
  {19.2, 25, 23.7},
  {18.7, 24.1, 23.6},
  {19, 23.2, 23.3},
  {18.1, 21.5, 22.9},
  {18, 20.6, 22.4},
  {16.9, 19.3, 21.1},
  {15.6, 18.2, 18.9},
  {15.1, 17.7, 17},
  {14.2, 17.3, 15.8},
  {14.2, 15.9, 15},
  {14.6, 16, 14.1},
  {13.9, 15.3, 13.5},
  {13.5, 15.4, 13},
  {14.2, 15.3, 12.7},
  {14.5, 15, 12.7},
  {14.6, 15.3, 13.2},
  {15, 15.7, 14},
  {15.9, 15.6, 15},
  {16.5, 16.2, 16.2},
  {16.7, 17.2, 17.8},
  {18, 18.4, 19.4},
  {18.5, 20.1, 21.6},
  {20, 20.8, 23.3},
  {20.5, 21.6, 23.4},
  {20.3, 21.1, 23.8},
  {18.2, 20.7, 23.4},
  {17.8, 19.3, 21.1},
  {17.1, 18.9, 20.1},
  {17.2, 18.3, 19.6},
  {15.6, 18, 18.9},
  {15.8, 17.5, 17.4},
  {16, 17.6, 16.4},
  {15.6, 17.3, 17},
  {15.5, 15.4, 17.2},
  {15.2, 15.2, 16.5},
  {15, 15.1, 15.9},
  {14.7, 14.4, 15.6},
  {14.5, 14.1, 15.4},
  {14.4, 14.2, 15.1},
  {14, 14.4, 14.9},
  {14, 14.4, 14.9},
  {14.2, 14.7, 15.9},
  {15, 15.9, 17.5},
  {16.4, 16.9, 19.3},
  {17, 18.6, 20.6},
  {18.6, 20.1, 21.3},
  {18.8, 20.9, 21.9},
  {18.8, 21.3, 22.1},
  {19, 21.4, 22.5},
  {18.9, 21.5, 22.1},
  {19, 21, 21.7},
  {18.4, 20.1, 22.1},
  {17.8, 19.4, 21.8},
  {17.3, 18.6, 20.9},
  {14.5, 17.7, 18.7},
  {14, 18, 17.1},
  {14.1, 17.8, 15.7},
  {15.3, 16.8, 15},
  {14.8, 17, 14.1},
  {13.3, 16.6, 13.6},
  {12.2, 14.8, 12.9},
  {11.4, 14.2, 12.3},
  {11.3, 13.4, 12},
  {10.9, 13.1, 11.8},
  {12.5, 13.1, 12.4},
  {13.4, 13.5, 13.7},
  {13.2, 14.8, 15.6},
  {13.3, 15.2, 17.3},
  {14.8, 15.4, 17.8},
  {15.6, 16, 18.1},
  {14.6, 16.1, 18},
  {14.2, 16, 18.5},
  {13.2, 16.5, 18.4},
  {13.9, 16.5, 17.9},
  {14.1, 16.5, 17.9},
  {14.2, 16.5, 17.9},
  {14.5, 15.9, 17.8},
  {14.3, 15.5, 18},
  {14.1, 14.8, 17.2},
  {13.7, 14.9, 15.8},
  {13.3, 14.7, 14.3},
  {12.5, 13.7, 13.2},
  {11.6, 13.3, 12.2},
  {10.7, 13.3, 11.2},
  {10.1, 13.3, 10.6},
  {10.2, 13.2, 10.3},
  {10.9, 13.1, 10.4},
  {11.4, 13.1, 10.5},
  {12.5, 13.6, 11.2},
  {13.6, 14.1, 12.4},
  {14.9, 14.6, 14.2},
  {16, 16, 16.4},
  {16.3, 16.9, 18},
  {14.9, 17.3, 18.2},
  {14.1, 16.9, 17.7},
  {14.7, 17.2, 18.4},
  {15.8, 17.5, 19.5},
  {16.8, 18.5, 19.9},
  {16.9, 18.6, 20.7},
  {16.3, 18.2, 20.3},
  {15.7, 17.5, 20},
  {14.9, 16.7, 18.9},
  {14.3, 16.2, 17.2},
  {14.3, 16, 15.3},
  {13.5, 15.3, 13.9},
  {12.3, 14.2, 12.7},
  {13.3, 13.3, 11.7},
  {11.5, 12.9, 11.1},
  {10.7, 12.7, 10.2},
  {10.1, 12.6, 9.8},
  {10, 12.5, 9.3},
  {11.4, 12.8, 9.4},
  {12.9, 13.9, 10.1},
  {14.2, 14.2, 12.4},
  {15.7, 15.7, 14.2},
  {16.8, 16.7, 17.6},
  {17.8, 18.6, 19.8},
  {18.9, 20.2, 21.5},
  {19.1, 21, 22.3},
  {18.7, 21.4, 22},
  {19.1, 22.2, 22.8},
  {18.7, 22.3, 23.3},
  {18.4, 22.5, 23.3},
  {18.3, 21.6, 22.7},
  {17.5, 20, 22.2},
  {16.2, 18.5, 20.4},
  {14.5, 17.7, 18.3},
  {14.1, 17.7, 16.6},
  {13.8, 17.7, 15.5},
  {13.1, 17.3, 14.6},
  {13.2, 16.8, 13.6},
  {12.5, 16.6, 12.9},
  {13.4, 16.3, 12.5},
  {13.7, 15.9, 12.1},
  {13.2, 15, 11.4},
  {13.7, 14.3, 10.9},
  {14.9, 15.5, 11.5},
  {15.2, 17.3, 15.2},
  {15.9, 19, 18.3},
  {16.5, 19.3, 20.8},
  {17.1, 20.3, 21.7},
  {16.6, 20.9, 21.7},
  {17, 20.3, 21.1},
  {17.1, 19.8, 21},
  {17.1, 19.7, 21.2},
  {17, 19.3, 20.8},
  {16.6, 19.2, 20.7},
  {14.8, 19, 20.2},
  {12.6, 17.4, 17.1},
  {12.5, 16.2, 14.7},
  {12.6, 15.5, 13.9},
  {12.6, 13.7, 13.6},
  {12.7, 13.6, 13.2},
  {11.9, 13.6, 13.1},
  {11.2, 13.2, 12.8},
  {10.6, 12.4, 12.3},
  {10.5, 11.9, 11.9},
  {10.9, 11.9, 11.5},
  {10.8, 11.6, 11.5},
  {10.7, 11.4, 11.8},
  {11, 11.4, 12.1},
  {10.8, 11.9, 12.6},
  {11.2, 12.3, 12.5},
  {12.3, 13.2, 12.4},
  {13.2, 13.6, 13.1},
  {13.6, 13.9, 14.1},
  {13.9, 15, 14.3},
  {12.8, 14.3, 13.5},
  {11, 11.1, 12.3},
  {10.4, 9.5, 12.7},
  {10.4, 11.4, 14.5},
  {10.3, 12.2, 15.4},
  {9.5, 11.9, 15.8},
  {7.8, 9.8, 12.9},
  {6.7, 8.7, 10.9},
  {6.4, 8.4, 9.5},
  {6.3, 8.9, 8.6},
  {6.4, 8.2, 8.2},
  {5.8, 7.6, 7.7},
  {5.5, 7.2, 7.2},
  {5.7, 7.4, 6.9},
  {5, 7.1, 6.9},
  {5.1, 7, 7},
  {5.9, 7, 7.5},
  {9.3, 7.2, 7.4},
  {10.5, 7.9, 7.8},
  {11.1, 10.7, 9.5},
  {12.3, 12.3, 13.1},
  {13.6, 14.2, 16.1},
  {14.7, 16.2, 17.6},
  {14.8, 17.2, 17.7},
  {14.2, 17, 18.2},
  {13.5, 16.3, 17.9},
  {13.9, 16.9, 18},
  {14.1, 17.5, 18.8},
  {14.2, 17, 18.2},
  {13.1, 15.6, 17.4},
  {12.2, 14.6, 16.5},
  {11.1, 13.3, 14.6},
  {10, 11.7, 12.4},
  {8.9, 11.3, 10.7},
  {8.6, 10.5, 9.8},
  {8.3, 9.8, 9},
  {8.3, 9.8, 8.4},
  {8.3, 10, 8.1},
  {8.1, 9.9, 7.7},
  {7.6, 9.4, 7.1},
  {9.1, 9.9, 7},
  {12.5, 9.5, 8.2},
  {13, 11.6, 11.1},
  {14.6, 15, 14.1},
  {16.6, 16.1, 17},
  {17.3, 17.3, 20.3},
  {18.2, 19.2, 22.9},
  {19.4, 21, 23.8},
  {20.1, 22.5, 23.6},
  {19.5, 22.1, 22.6},
  {18.8, 21.9, 22.9},
  {18.2, 20.8, 23.3},
  {17.2, 20.5, 22.3},
  {16.5, 19.6, 21.4},
  {16, 18.2, 20.1},
  {14.5, 16.6, 17.7},
  {14.1, 16, 15.5},
  {13.3, 16, 14.2},
  {12.7, 15.8, 13.4},
  {12.8, 15.6, 12.6},
  {12, 14.5, 11.9},
  {11.9, 13.9, 11.6},
  {12.1, 14.1, 11.2},
  {12, 13.7, 10.9},
  {12.8, 14.3, 10.4},
  {14.2, 14.3, 11},
  {16, 14.7, 12.7},
  {17.3, 15.7, 14.7},
  {17.5, 17.7, 16.4},
  {19.1, 18.9, 18.6},
  {20.2, 19.3, 21.2},
  {19.9, 21, 23},
  {20.5, 24.2, 24.3},
  {22, 24.4, 26.6},
  {22.6, 25.7, 27.2},
  {22.1, 25.5, 25.9},
  {20.8, 25, 25.1},
  {19.5, 22.8, 23.5},
  {16.7, 20.5, 21.2},
  {15.8, 18.4, 18.5},
  {15.4, 17.3, 16.4},
  {14.1, 16.8, 15},
  {13.1, 15.8, 14.1},
  {12.6, 14.7, 13.2},
  {12, 14.2, 12.3},
  {11.7, 13.5, 11.6},
  {11.4, 12.8, 11},
  {11.5, 12.8, 10.6},
  {12.4, 13.2, 10.3},
  {16.3, 13.5, 11.2},
  {17.3, 15, 13.9},
  {17.6, 16.2, 16.5},
  {18.4, 17.5, 18.6},
  {19.7, 19.3, 21.5},
  {20.5, 21, 23.4},
  {21.9, 22.3, 24.5},
  {21.7, 22.9, 24.2},
  {21.4, 22.6, 23.6},
  {21.4, 22.4, 23.7},
  {20.3, 21.9, 23},
  {19.2, 22.1, 23.2},
  {19.3, 21.2, 23.1},
  {18.4, 19.2, 20.5},
  {17.7, 17.5, 18.2},
  {15.4, 17.7, 16.3},
  {13.6, 17.8, 15},
  {13.7, 17.3, 14.2},
  {13.2, 16.9, 13.4},
  {12.8, 16.2, 12.8},
  {13.2, 16.1, 12.6},
  {12.9, 15.6, 12.6},
  {12.7, 15.2, 12.6},
  {13.8, 15.2, 12.6},
  {14.3, 15.3, 13},
  {14.9, 15.5, 14},
  {14.9, 15.7, 15.2},
  {15.5, 15.6, 16.6},
  {15, 15.5, 17.7},
  {14.5, 15.9, 19.5},
  {14.2, 15, 18.7},
  {13.6, 12.8, 15.8},
  {13.2, 11.1, 14.7},
  {12.1, 12.7, 13.9},
  {12.5, 12.4, 15.2},
  {12.4, 11.5, 15.3},
  {12.1, 12.3, 14.7},
  {11.5, 10.8, 14.5},
  {11.2, 9.9, 14.2},
  {10.9, 9.8, 13.6},
  {10.9, 9.8, 13},
  {10.4, 9.8, 12.5},
  {9.8, 9.8, 11.8},
  {9, 9.6, 11.5},
  {7.8, 9.2, 11},
  {7.8, 8.5, 11.1},
  {7.6, 8.2, 10.9},
  {6.9, 7.8, 9.9},
  {7.1, 8.5, 10},
  {7.4, 9.2, 11},
  {7.3, 9.2, 11.4},
  {8, 10, 11.6},
  {9, 11.6, 13.7},
  {9.6, 12.5, 14.2},
  {8.4, 12.1, 12.7},
  {6.5, 12.8, 11.9},
  {5.2, 12.4, 10.3},
  {6.5, 12.3, 10.6},
  {7.4, 12.1, 10.8},
  {7.2, 11.4, 11.3},
  {7.3, 10.9, 11.2},
  {5.3, 9.4, 10.3},
  {3.9, 8, 8},
  {4.2, 7.7, 6},
  {4.2, 7.3, 4.7},
  {3.1, 6.6, 3.8},
  {2.6, 6.4, 2.9},
  {1.6, 5, 2.3},
  {1.3, 4.3, 1.5},
  {1.6, 4.2, 1},
  {2, 3.7, 0.6},
  {3.9, 3.9, 0.4},
  {5.9, 4, 1},
  {7.3, 5.9, 4},
  {8.5, 9.5, 7.7},
  {10.9, 11.3, 11.5},
  {11.2, 12.9, 14.4},
  {10.2, 14.2, 15.6},
  {9.1, 13.6, 13.8},
  {8.5, 13.5, 14},
  {8.6, 12.9, 15.1},
  {10.7, 12.4, 15.3},
  {10.7, 12.3, 14.3},
  {10.2, 12.1, 14.4},
  {8.3, 11.4, 13.3},
  {6.6, 9.4, 12.2},
  {5.4, 7.9, 10.7},
  {5, 6.8, 8.7},
  {5.1, 6.9, 7.2},
  {6.2, 7.3, 5.8},
  {5.9, 7, 5.2},
  {4.5, 6.3, 4.4},
  {4.9, 5.3, 3.5},
  {4.9, 5, 2.6},
  {3.2, 4.8, 2.1},
  {5.2, 5.2, 1.5},
  {7.3, 6.4, 2.6},
  {7.9, 7.7, 6.6},
  {9.9, 10.6, 10.6},
  {11.8, 12.7, 13.7},
  {11.8, 14.3, 15.6},
  {13.4, 15.4, 17},
  {14.2, 16.6, 17.9},
  {14.4, 16.8, 19},
  {13.6, 17.6, 19.2},
  {13.2, 16.5, 18.1},
  {11.7, 14.9, 16.4},
  {11.1, 12.4, 15.1},
  {9.5, 10.4, 12.3},
  {5.9, 10.1, 9.3},
  {4.4, 8.6, 7.8},
  {3.7, 7.5, 7.4},
  {3.3, 6.2, 7.2},
  {3.3, 5.7, 7},
  {3.9, 5, 6.9},
  {4.2, 5.2, 6.6},
  {4.7, 5.5, 6.3},
  {4.6, 5.8, 6},
  {4.9, 6.3, 5.9},
  {4.8, 6.9, 5.9},
  {5.9, 8.3, 6.4},
  {8.5, 9, 7.4},
  {9.9, 10.7, 9.5},
  {11.5, 12.2, 12},
  {12.7, 13.6, 15.5},
  {13.5, 14.7, 16.5},
  {13.7, 15.4, 17.5},
  {13.2, 16.1, 18.2},
  {12.5, 16.7, 18.6},
  {14.5, 16.1, 18.8},
  {13.7, 14.9, 18},
  {12.5, 13.3, 16.7},
  {10.7, 12.1, 15.8},
  {10.5, 11.4, 15.1},
  {10.3, 10.8, 14.7},
  {10.1, 10.7, 14},
  {9.9, 10.3, 13.8},
  {10, 10.3, 13.6},
  {10.1, 10.2, 12.4},
  {10.3, 10.2, 11.1},
  {10.6, 10.2, 10.4},
  {10.6, 10.1, 9.7},
  {10.8, 9.8, 9},
  {10.5, 10.1, 10.7},
  {10.2, 10.5, 12.4},
  {10.4, 11.2, 12.8},
  {11.4, 12.7, 14.2},
  {12.3, 13.3, 15.1},
  {12.4, 14.2, 16.4},
  {13.5, 14.5, 17.3},
  {14.1, 14.8, 17.6},
  {14.2, 15, 18.3},
  {13.5, 15.2, 17.9},
  {14.1, 15.3, 18},
  {14.2, 15.3, 18.5},
  {13.5, 15.8, 18},
  {12.8, 14.6, 17.6},
  {12.2, 13.9, 17.2},
  {11.4, 12.6, 16.6},
  {10.2, 11.7, 15.1},
  {8.5, 11.3, 13},
  {7.1, 11.1, 10.1},
  {7.9, 10.7, 8.4},
  {7.4, 10.2, 7.4},
  {6.1, 9.3, 6.6},
  {6.2, 9.5, 5.7},
  {6.5, 10.1, 5.8},
  {7.8, 9.9, 6.1},
  {8.4, 10.3, 6.9},
  {10.3, 10.5, 8.3},
  {11.9, 11.7, 10.5},
  {12.7, 14.1, 13.3},
  {14.3, 16, 16.2},
  {15.7, 17.7, 19.1},
  {16.7, 18.7, 20.7},
  {17.2, 19.6, 21.5},
  {16.6, 19.5, 21.8},
  {15.7, 19.8, 20.4},
  {16.2, 20.3, 21},
  {15.5, 19.8, 21.5},
  {14.6, 18.2, 19.3},
  {13.2, 16.2, 17.8},
  {11.6, 14.7, 15.8},
  {10.9, 14, 13.1},
  {11.2, 13.6, 11.4},
  {9.7, 13.5, 10.4},
  {9.9, 13.1, 9.9},
  {9.8, 12.5, 9.6},
  {9.4, 11.8, 9.1},
  {8.9, 11.8, 8.9},
  {8, 11.5, 8.7},
  {8.4, 11.6, 8.4},
  {10.9, 11.7, 9.5},
  {12.7, 12.6, 11.5},
  {13.2, 14, 13.1},
  {14.1, 15.7, 15.1},
  {15.8, 16.7, 18.1},
  {16.5, 17.5, 19.8},
  {15.4, 18, 21.2},
  {16, 18.4, 20.3},
  {15.6, 18.9, 19.6},
  {14.6, 19.4, 19.9},
  {13.9, 17.4, 18.8},
  {13.2, 15.4, 16.8},
  {12.6, 15, 16.2},
  {10.6, 13.7, 15.9},
  {8.9, 13, 14.6},
  {8.7, 12.7, 13.1},
  {8.3, 12.2, 12},
  {7.3, 11.3, 10.7},
  {7.1, 10.2, 9.5},
  {6.7, 9.5, 8.4},
  {6.8, 8.7, 7.7},
  {6.5, 8.1, 7.7},
  {6.1, 7.8, 7.8},
  {7.3, 8.2, 8},
  {9.8, 9.9, 9.3},
  {9.6, 10.2, 10.8},
  {10.3, 11.1, 12.7},
  {11.9, 12.8, 15.4},
  {12.6, 14.7, 17.3},
  {14.2, 16.3, 18.2},
  {13.8, 16.7, 17.4},
  {14, 18.1, 19.1},
  {14.5, 18.1, 19.9},
  {14.8, 17.7, 18.8},
  {14.7, 16.8, 18.7},
  {13.4, 15.4, 18.1},
  {12.5, 14.3, 17.6},
  {11.3, 13.5, 16.5},
  {10.2, 12.6, 15.5},
  {8.7, 12, 14.9},
  {8.2, 11.1, 14},
  {7.6, 9.7, 13.7},
  {4.7, 8.5, 13},
  {5.1, 7.4, 11.5},
  {4.8, 7.1, 9.6},
  {4.4, 7.1, 8.1},
  {3.8, 5.9, 7},
  {4.8, 6.6, 6.3},
  {7.7, 6.9, 6.9},
  {10.1, 9.4, 10.4},
  {10.7, 12.6, 12.8},
  {11.8, 14.7, 16.2},
  {13.3, 16.1, 17.3},
  {14, 17.7, 18.7},
  {13.9, 19, 19.6},
  {13.7, 19.6, 19.2},
  {14.4, 20.1, 18.9},
  {14.1, 18.3, 18.9},
  {13.8, 17.4, 18.3},
  {13.3, 16.6, 18.1},
  {12, 15.6, 17.2},
  {11.2, 13.8, 16},
  {10.6, 12.5, 14.6},
  {9.6, 11.4, 12.6},
  {8.3, 10.8, 11},
  {7.6, 10.9, 10.2},
  {7.1, 10.3, 9.6},
  {7.4, 9.2, 8.5},
  {7.4, 8.2, 8},
  {7.9, 8.2, 7.8},
  {8.2, 8.6, 7.6},
  {9.1, 8.9, 7.8},
  {10.9, 8.9, 9.8},
  {10.9, 10.4, 12},
  {12, 14, 13.8},
  {13.3, 15, 16.6},
  {14.1, 16.2, 18.4},
  {14.8, 17.9, 18.8},
  {15.4, 19.2, 19.9},
  {16.2, 19.9, 20.9},
  {15.9, 19.8, 21.1},
  {15.7, 19.5, 20.2},
  {15.4, 18.6, 19.9},
  {14.3, 17.1, 19.3},
  {13.3, 16.1, 18.2},
  {13, 15.1, 17.6},
  {12.7, 13.9, 17.2},
  {12.1, 13.4, 16.5},
  {11.7, 13.3, 16.1},
  {11.4, 13.3, 15.7},
  {11.2, 13.3, 15.2},
  {10.5, 12.9, 14.6},
  {9.8, 12.4, 14.3},
  {9, 10.2, 13.8},
  {9, 9.5, 13.6},
  {9, 9.6, 13.5},
  {10.9, 10.2, 13.6},
  {12.5, 11.2, 14.7},
  {13.2, 13.7, 16.5},
  {14.3, 15.3, 16.8},
  {14.2, 16, 17.8},
  {14.5, 17.7, 19.3},
  {14.6, 18.7, 19.7},
  {15.9, 18.9, 20.2},
  {16, 19.1, 20},
  {15.9, 19, 19.5},
  {15.4, 18.5, 19.5},
  {14.3, 17.6, 19.1},
  {13.2, 16.5, 18.5},
  {12.3, 14.9, 17.6},
  {11.3, 13.8, 15.7},
  {9.7, 13, 13.8},
  {9.9, 12.3, 12.9},
  {8.8, 12.2, 12.1},
  {8.6, 12.3, 10.7},
  {8.9, 10.6, 10.5},
  {8.7, 9.5, 9.9},
  {8.3, 9.5, 8.8},
  {8, 9.6, 7.8},
  {8.9, 9.9, 7.6},
  {11.8, 10.8, 8.8},
  {12.5, 12.1, 12.5},
  {13.3, 14.1, 15},
  {14.6, 15.5, 16.6},
  {16.5, 16.3, 18},
  {17.8, 18.2, 20.1},
  {18.6, 20.2, 21.9},
  {19.8, 22, 23.9},
  {19.9, 23.5, 25.4},
  {19.3, 24.8, 25.3},
  {18.8, 25, 23.8},
  {17.3, 23.9, 23.7},
  {16.5, 20.5, 23.3},
  {14.6, 19.4, 21.6},
  {14, 18.3, 19.7},
  {13.6, 17.5, 18},
  {13, 16.7, 16.4},
  {12.7, 15.8, 14.8},
  {13.2, 15.7, 13.6},
  {12.6, 14.9, 12.8},
  {12.3, 14.2, 11.7},
  {11.7, 13.6, 11.6},
  {10.9, 13.1, 11.9},
  {11.5, 12.5, 12},
  {11.9, 13.3, 12.8},
  {13, 14.6, 15},
  {13.8, 16.2, 17.7},
  {14, 17.7, 18.3},
  {15, 18.3, 19},
  {15, 19, 19.7},
  {15.5, 19.4, 19.8},
  {15.6, 19.8, 20.4},
  {16.1, 20, 20.7},
  {16.4, 19.9, 20.6},
  {15.6, 19.2, 20.4},
  {14.9, 18.2, 19.6},
  {14.2, 17.3, 18.9},
  {13.7, 16.2, 18.4},
  {13.3, 15.2, 18},
  {13.4, 14.8, 17.6},
  {12.9, 15, 16.2},
  {12.3, 14.9, 15},
  {11.4, 14.4, 14.7},
  {10.5, 14, 14.1},
  {10.1, 12.8, 13.3},
  {9.5, 12.6, 12.5},
  {9.5, 11.6, 12.2},
  {10.6, 11.5, 11.3},
  {13.4, 12.3, 12.2},
  {14.4, 13.8, 15.2},
  {14.7, 16.1, 17.4},
  {15.5, 17.2, 19.6},
  {17.3, 18.9, 22},
  {17.9, 20.9, 23.4},
  {19, 22.1, 23.5},
  {19.7, 22.6, 24},
  {19.9, 22.8, 23.8},
  {19.3, 22.5, 23.2},
  {18.4, 21.8, 23.1},
  {17.6, 21, 22.7},
  {16.4, 20, 22.2},
  {15.9, 18.5, 21.2},
  {15.5, 17.1, 19.7},
  {14.8, 16.3, 17.1},
  {13.3, 15.4, 15.1},
  {12.2, 14.9, 13.9},
  {11.4, 14.5, 12.9},
  {11, 14.1, 12.1},
  {10.9, 13.1, 11.5},
  {10.7, 12.2, 10.9},
  {10.7, 12.1, 10.4},
  {12.1, 12.8, 10.2},
  {15.6, 13.6, 11.6},
  {16.6, 16, 14.5},
  {16.8, 18, 17.1},
  {18.6, 20, 20.2},
  {20, 20.7, 23.1},
  {21.2, 23, 25.2},
  {22.4, 25, 26.5},
  {22.7, 25.4, 25.7},
  {22.4, 25.3, 26.2},
  {20.1, 24.6, 26},
  {19.2, 22.9, 22.5},
  {18.5, 22.6, 20.1},
  {18.4, 21.8, 18.8},
  {17.7, 19.9, 18.5},
  {15.1, 18.7, 17.3},
  {16.6, 18.1, 16.1},
  {14.7, 17.7, 15.7},
  {14.1, 17.2, 14.8},
  {13.9, 16.6, 14.1},
  {13.1, 16.1, 13.4},
  {12.9, 14.9, 12.8},
  {12.7, 14.5, 12.2},
  {12, 14.1, 11.6},
  {13.4, 14.7, 11.5},
  {17.4, 15.1, 12.7},
  {18.7, 16.3, 14},
  {19.7, 18.2, 16.6},
  {20.6, 20.4, 19.9},
  {21.5, 22.2, 23.2},
  {22.4, 24.2, 25.7},
  {23.2, 26.3, 27.4},
  {23.3, 26.8, 26.9},
  {22.8, 26.3, 27},
  {22.8, 25.8, 26.9},
  {22.9, 25.5, 26.9},
  {21.7, 24.7, 27.1},
  {20.3, 23.5, 26.1},
  {19.8, 21.9, 24.4},
  {19.4, 20.5, 22.3},
  {18.1, 19.7, 19.6},
  {15.9, 19.7, 18.3},
  {15.4, 18.7, 17},
  {15.1, 18, 15.8},
  {14.7, 17.6, 15.2},
  {14.6, 16.3, 14.4},
  {14, 16.1, 13.9},
  {13.7, 15.8, 13.3},
  {15.1, 16, 13},
  {18.9, 16.4, 14.1},
  {20, 18, 17.6},
  {20, 19.8, 20.5},
  {20.8, 21.4, 22.9},
  {21.8, 23.4, 25.3},
  {23.3, 25.3, 26.8},
  {23.5, 26, 26.8},
  {23.8, 26.4, 27},
  {24.5, 26.7, 27.5},
  {23.6, 26.4, 27.7},
  {22.3, 25.4, 27.5},
  {21.6, 24.7, 27.2},
  {20.5, 23.9, 26.3},
  {19.8, 22.4, 24.8},
  {18.4, 21.1, 22.4},
  {17.1, 20.4, 19.6},
  {15.8, 19.8, 18},
  {14.9, 19.3, 16.6},
  {14.5, 18.6, 15.6},
  {14.8, 17.9, 14.7},
  {14.8, 17.6, 14},
  {14, 17, 13.3},
  {13.9, 16, 12.6},
  {16.1, 16.1, 12.7},
  {18.1, 17.4, 14.7},
  {19.9, 18.5, 17.2},
  {20.4, 20.2, 20},
  {20.6, 21.5, 21.7},
  {21.9, 22.9, 24.5},
  {22.6, 24.6, 26.6},
  {22.9, 25, 26.8},
  {22.2, 25.3, 27.4},
  {22.8, 24.2, 25.8},
  {21.9, 25.2, 26.7},
  {22.3, 24.7, 26.4},
  {21.6, 24.2, 26},
  {20.3, 23.1, 25},
  {18.5, 22, 23.8},
  {17, 20.9, 22.8},
  {16.2, 19.4, 20.6},
  {15.9, 18.4, 17.7},
  {15, 18.4, 16.7},
  {14.1, 17.8, 15.2},
  {13.4, 17.4, 14.3},
  {13.2, 16.5, 13.6},
  {13.2, 15.6, 12.9},
  {12.9, 15.2, 12.2},
  {14.4, 15.5, 12.1},
  {17.6, 16.1, 13.4},
  {18.3, 17.4, 16.4},
  {20.1, 19.2, 19.2},
  {20.6, 20.1, 22.1},
  {21.6, 22.2, 24.3},
  {22.9, 23.9, 26.3},
  {23.5, 25.9, 27},
  {23.2, 25.7, 26.9},
  {23.6, 25.8, 27.5},
  {22.8, 24.8, 27.4},
  {22.9, 24.7, 27.9},
  {22.5, 21.3, 27.1},
  {21, 21.5, 26.6},
  {19.6, 20.7, 24.7},
  {18.6, 19.7, 23},
  {17.9, 19.6, 21.3},
  {16.9, 18.4, 19.2},
  {16.3, 18.1, 18},
  {15.1, 17.5, 17},
  {14.8, 17.2, 16.2},
  {14.6, 16.5, 15.9},
  {14.1, 16.2, 14.7},
  {14, 15.7, 14.2},
  {16.2, 15.9, 14},
  {19.2, 16.3, 15.1},
  {19.8, 17.4, 18.6},
  {19.7, 19.1, 21.8},
  {21.4, 21.6, 24},
  {22.1, 23.7, 25.8},
  {22.7, 24.5, 25.6},
  {24.3, 25.4, 27.6},
  {23.4, 27.5, 28.4},
  {23.8, 25.5, 26.3},
  {24, 23.6, 27.2},
  {23.3, 24.8, 27.7},
  {21.6, 24.7, 26.6},
  {20.7, 24, 26.4},
  {19.6, 22.5, 25.2},
  {18.1, 20.7, 23.5},
  {17, 20.4, 20.9},
  {16.5, 19.4, 19.4},
  {16, 18.6, 18.3},
  {15.6, 17.9, 17.3},
  {15.2, 17.9, 16.5},
  {14.7, 17.1, 15.8},
  {14.4, 16.4, 15.2},
  {14.7, 16.1, 14.6},
  {15.7, 16.3, 14.5},
  {19.3, 16.9, 15.7},
  {20.6, 18.1, 18.8},
  {21.9, 20.6, 21},
  {22.4, 21.9, 24.1},
  {23.2, 24, 26.3},
  {23.7, 25.5, 26.2},
  {24.2, 26.6, 27.5},
  {23.7, 27.3, 27.9},
  {23.2, 26.8, 27.4},
  {23.7, 26.4, 27.2},
  {22.6, 26, 27.2},
  {22.5, 25.2, 26.4},
  {21.6, 24.4, 26},
  {20.6, 23.3, 25.9},
  {20.1, 22.3, 23.9},
  {19.8, 20.7, 21.3},
  {19.5, 20.4, 19.2},
  {19.2, 20.9, 18},
  {17.2, 19.6, 17.3},
  {15.8, 19.5, 16.5},
  {15.7, 18.8, 16},
  {16.2, 18.1, 15.5},
  {15.7, 17.5, 14.9},
  {16.1, 17.4, 14.9},
  {19.8, 18, 16},
  {20.8, 19.2, 19},
  {21.3, 21.2, 21},
  {22.4, 22.4, 24.2},
  {23.3, 23.9, 26.6},
  {24.7, 25.6, 28.2},
  {25.4, 27.4, 29.2},
  {26.4, 28, 29.5},
  {26.7, 27.8, 29.7},
  {25.3, 26.9, 29.2},
  {23.9, 25.8, 28.5},
  {23.1, 25.4, 27.9},
  {22.8, 24.8, 27},
  {22.5, 23.4, 26.2},
  {20.3, 22.4, 24.4},
  {18.8, 22.3, 22.9},
  {18.2, 22, 21.3},
  {17.4, 21.5, 20.2},
  {17.2, 21.4, 19},
  {17.3, 20.9, 18.2},
  {16.9, 20, 17.4},
  {17.4, 19, 16.9},
  {17.6, 18.3, 16.5},
  {18.2, 18.8, 16.2},
  {20.1, 20, 17.3},
  {21.3, 20.6, 19.6},
  {21.8, 21.7, 21.6},
  {22.4, 22.5, 23},
  {23, 23.5, 25.2},
  {24.5, 25, 27.3},
  {25.3, 26.5, 28.5},
  {26.1, 28.1, 30.2},
  {25.7, 27.6, 29.1},
  {24.9, 28, 29.8},
  {25.5, 27.7, 29.5},
  {24.8, 27.1, 29.1},
  {23.2, 26, 28.4},
  {22.3, 25, 27.6},
  {21.7, 24.2, 25.5},
  {21.2, 23.5, 22.2},
  {20.7, 22.6, 20.2},
  {20.1, 21.3, 18.8},
  {19, 21.1, 17.9},
  {17.7, 20.9, 17},
  {16.6, 20.1, 16.4},
  {16.4, 19.3, 16},
  {16.5, 18.6, 15.4},
  {17.7, 18.3, 15.2},
  {20.4, 19, 16.3},
  {21.7, 20, 19.6},
  {22.6, 22.2, 22.2},
  {23.4, 23.5, 24.9},
  {23.4, 25.5, 27.6},
  {24.3, 25.7, 25.6},
  {24.2, 25.7, 25.1},
  {24.9, 27.1, 26.4},
  {23.1, 25.5, 20.8},
  {22.5, 25, 19.7},
  {23.3, 25.5, 22.2},
  {23.9, 26.1, 24.5},
  {22, 24.4, 21.6},
  {21.6, 23.3, 20.6},
  {19.3, 22, 19.4},
  {18.7, 20.6, 18.6},
  {18.8, 20.3, 18.3},
  {19.2, 20.3, 17.9},
  {19.3, 19.9, 17.5},
  {18.9, 19.2, 17.1},
  {17.7, 18.4, 16.7},
  {17.3, 18.3, 16.1},
  {17.2, 17.9, 15.5},
  {18.1, 17.9, 15.2},
  {19.2, 18.9, 16.1},
  {19.7, 20.5, 19.2},
  {20.1, 22.7, 21.2},
  {21.5, 23.5, 23.1},
  {23.1, 24.3, 25.6},
  {24.7, 26.1, 27.7},
  {25.1, 27.3, 28.5},
  {25.5, 27.6, 28.1},
  {25, 28.1, 28.1},
  {24.4, 27.9, 27.9},
  {24.6, 27.7, 28.1},
  {24.2, 26.9, 27},
  {23, 25.8, 26.6},
  {21.9, 24.1, 25.3},
  {19.2, 22.9, 21.5},
  {18.7, 22.8, 19.6},
  {18.7, 22.3, 18.5},
  {18.3, 21.6, 17.4},
  {18.8, 21.4, 16.5},
  {19, 21.4, 16.3},
  {19.6, 21.4, 17},
  {18.8, 20.3, 17.2},
  {17.1, 19, 16.4},
  {17.3, 18.8, 15.6},
  {20.9, 19.3, 16.6},
  {21.9, 20.3, 19.9},
  {22.8, 22.9, 22.6},
  {23.9, 24, 25.1},
  {25.1, 25.8, 27.3},
  {25.4, 27.4, 28.9},
  {26, 28.4, 28.9},
  {25.6, 28.8, 29.3},
  {25.8, 28.8, 29.5},
  {25.5, 29, 28.5},
  {25.3, 28.4, 28.7},
  {24.9, 27.4, 28.3},
  {23.5, 26.3, 27.3},
  {22.5, 24.9, 26.6},
  {22.1, 24, 24.3},
  {21.4, 22.9, 22.4},
  {19.7, 22.7, 20.5},
  {19, 22.5, 19.9},
  {15.9, 19.5, 19.8},
  {15.5, 18.1, 19.1},
  {15.6, 17.7, 18.2},
  {15.9, 17.4, 17.8},
  {15.3, 17, 17.8},
  {15.1, 16.9, 17.7},
  {15.1, 16.8, 17.8},
  {16.4, 17.3, 17.9},
  {18.1, 18.4, 19},
  {20.4, 20.2, 21.3},
  {21.7, 21.8, 24.1},
  {23.6, 23.3, 25.7},
  {23.6, 24.8, 27.6},
  {25.3, 26.6, 29},
  {25.5, 27.7, 29.2},
  {22.9, 27, 28},
  {22.5, 25.1, 26},
  {23.7, 25.4, 26.4},
  {21.9, 24.8, 26.9},
  {20.9, 22.6, 24.8},
  {18.6, 21.1, 22.2},
  {18.2, 20.2, 20.4},
  {19.2, 19.3, 19.4},
  {18.8, 19.2, 19.3},
  {19, 18.9, 18.9},
  {19.3, 18.6, 18.7},
  {19.2, 17.7, 18},
  {18.7, 17.1, 17.4},
  {18.8, 17, 16.7},
  {19.5, 17.2, 16.3},
  {21.3, 17.7, 17.5},
  {23, 18.9, 20},
  {23.7, 21.6, 22.7},
  {24.7, 23.5, 25},
  {24.4, 24.8, 27.8},
  {25.3, 26.9, 29.6},
  {25.6, 28.5, 29.9},
  {25.7, 29.2, 30.2},
  {25.4, 29.1, 30},
  {25.6, 28.6, 29.7},
  {25.4, 28.1, 29.7},
  {24.9, 27.8, 29},
  {23.6, 26.7, 28.1},
  {22.4, 24.9, 26.1},
  {19.5, 23, 22.2},
  {20.2, 22.7, 20.2},
  {18.9, 22.2, 18.8},
  {17.8, 20.9, 17.5},
  {18.2, 20, 16.8},
  {17.1, 19.1, 16.1},
  {16.6, 18, 15.4},
  {16.8, 17.5, 14.7},
  {16.2, 17.5, 14.2},
  {17.5, 17.9, 14},
  {20.7, 18.3, 15.1},
  {22.1, 19.3, 18.7},
  {22.9, 21.5, 21.8},
  {24.8, 24, 24.4},
  {25.1, 26.3, 27.1},
  {26, 27.8, 29.4},
  {26.4, 28.9, 30.2},
  {25.9, 29.2, 30.4},
  {25.6, 29, 30.3},
  {25.6, 29.1, 30.4},
  {25.7, 28.7, 30.1},
  {24.9, 27.6, 29.4},
  {23.9, 26.5, 29.1},
  {23.1, 25.7, 28},
  {21.8, 24.3, 25.7},
  {20.9, 23.2, 22.2},
  {20.7, 22.8, 20.5},
  {18.5, 21.5, 20.1},
  {18.8, 21, 18.9},
  {19.3, 20.8, 18.7},
  {19.1, 19.8, 18.1},
  {18.6, 19.6, 17.3},
  {19.2, 20, 17.1},
  {19.2, 17.6, 17.7},
  {18.8, 16.8, 17.8},
  {19.9, 17.1, 18.5},
  {19.7, 18.5, 19.6},
  {20.6, 20.5, 22.2},
  {22.1, 20.7, 24.5},
  {23.3, 22.5, 26.6},
  {24.4, 24.9, 28.3},
  {25.3, 26, 29.8},
  {26, 26.5, 30.3},
  {26.4, 27.5, 30.3},
  {25.1, 27.9, 29.3},
  {24, 27.6, 28.6},
  {23, 26.3, 27.9},
  {22.1, 24.9, 27.2},
  {22.2, 23.8, 25.1},
  {21.2, 23.1, 22.3},
  {19.3, 22.7, 20.9},
  {18.4, 21.4, 19.9},
  {18.3, 20.1, 19.1},
  {19.2, 20.2, 18.6},
  {19, 20.7, 19.3},
  {18.2, 19.9, 19.2},
  {15.9, 19.9, 18.5},
  {15.9, 18.4, 18.6},
  {16.1, 17.1, 18.3},
  {16.1, 15.1, 18.2},
  {15.5, 14.3, 17.8},
  {14.9, 14.3, 17.2},
  {14.9, 14.5, 16.7},
  {13.8, 14.4, 16.8},
  {13.6, 14.3, 16.7},
  {14.7, 14.4, 16.6},
  {15.9, 16.1, 18.5},
  {16.6, 17.7, 21.7},
  {17.9, 17.8, 23.5},
  {18.4, 18.6, 23.5},
  {16, 18.3, 23.4},
  {15.3, 17.3, 21.1},
  {15.7, 15.8, 18.2},
  {14.5, 15.7, 16.4},
  {14.4, 15.5, 15.3},
  {13.4, 15.1, 14.5},
  {13.8, 14.3, 13.7},
  {12.7, 13.5, 13},
  {11.9, 13.6, 12.3},
  {12.2, 13.7, 11.9},
  {11.9, 13.4, 11.4},
  {14.2, 13.4, 11.1},
  {16.8, 13.8, 11.8},
  {17.4, 15.2, 14.3},
  {18.2, 17.8, 17.9},
  {19.5, 20.7, 21.2},
  {21.1, 22.6, 24.5},
  {22.8, 24.6, 26.7},
  {23.8, 25.5, 27.6},
  {24.7, 26.8, 28.4},
  {25.2, 27.6, 29.5},
  {25.8, 28.1, 30.5},
  {25.7, 28.1, 30.2},
  {23.3, 27.9, 28.2},
  {21.7, 25.1, 25.9},
  {20.9, 22.9, 25.3},
  {18.9, 21.6, 21.9},
  {18.4, 20.6, 21.1},
  {17.6, 20.8, 19.3},
  {17.8, 20, 17.5},
  {16.3, 19, 16.5},
  {16.4, 18.4, 15.5},
  {15.8, 17.7, 14.7},
  {15.2, 17.4, 13.8},
  {15.2, 17, 13.3},
  {16.3, 16.5, 12.8},
  {19.1, 16.9, 14},
  {19.3, 18, 17.3},
  {19.8, 20.9, 20},
  {21, 22.8, 22.7},
  {22.1, 23.8, 25.3},
  {22.9, 25.1, 27},
  {23.4, 25.9, 27.1},
  {23.3, 26.9, 27.3},
  {22.6, 26.4, 27.7},
  {22.7, 26.5, 27},
  {21.9, 25.5, 26.6},
  {21.7, 24.4, 25.9},
  {21.3, 23.7, 26.1},
  {20.2, 22.6, 25.2},
  {19, 21.7, 23},
  {18.7, 20.4, 21.1},
  {17.3, 20.5, 20.3},
  {17, 20.7, 19.5},
  {16.8, 19.9, 18.8},
  {16.9, 19.7, 18.8},
  {16.6, 19, 19.1},
  {16.7, 17.7, 18.9},
  {16.8, 17.4, 19},
  {16.8, 17.8, 19.1},
  {17.3, 18.6, 19.5},
  {18.5, 19.1, 20.5},
  {18.8, 20.6, 22.2},
  {20, 21.7, 23.7},
  {20.7, 22.7, 24.4},
  {21.2, 24.1, 25},
  {21.8, 24.7, 25.1},
  {22.2, 25, 25.3},
  {21.7, 25, 25.5},
  {21.4, 24.9, 25.4},
  {19.9, 24.3, 25.2},
  {19.2, 22.9, 23.8},
  {18.9, 22.1, 23.2},
  {18.6, 20.9, 22.5},
  {17.2, 19.4, 20.4},
  {16.7, 19.7, 19.3},
  {16.9, 19.8, 18.8},
  {16.9, 17.7, 18.5},
  {16.3, 17.5, 18.3},
  {15.5, 17.8, 17.8},
  {15.2, 17.9, 16.8},
  {14.3, 17.4, 15.8},
  {15.1, 17, 15.2},
  {15.1, 17.3, 15.3},
  {17.5, 18.4, 16.4},
  {18.3, 19.1, 18.1},
  {19, 20.5, 19.7},
  {19.8, 21.4, 22},
  {20.5, 23, 24.4},
  {21.3, 24, 25.8},
  {22, 24.9, 26.2},
  {22.9, 25.5, 26.8},
  {22.3, 25.8, 26.7},
  {21.7, _, 26.1},
  {20, _, 24},
  {20.5, _, 24.7},
  {19.9, _, 24.1},
  {18.6, _, 21.6},
  {16.9, _, 19.6},
  {16.6, _, 19.2},
  {16.4, _, 17.7},
  {15.5, _, 17.3},
  {14.5, _, 16.9},
  {14.1, _, 15.9},
  {14.1, _, 15.1},
  {13.9, _, 14.9},
  {14, _, 15.2},
  {13.8, _, 15.1},
  {15.3, _, 15.2},
  {17.1, _, 15.5},
  {19, _, 16.4},
  {19.6, _, 18.8},
  {20.4, _, 21.8},
  {21.1, _, 24.4},
  {21.9, _, 25.8},
  {22.3, _, 25.7},
  {22.5, _, 25.1},
  {21.7, _, 25.1},
  {21.1, _, 24.7},
  {19.9, _, 23.9},
  {19.5, _, 24.1},
  {19.1, _, 22.4},
  {18, _, 21.6},
  {17.5, _, 21.7},
  {16.6, _, 21.6},
  {17.2, _, 20.6},
  {17, _, 20.2},
  {16.5, _, 19.5},
  {16.5, _, 19},
  {16.7, _, 18.9},
  {16, _, 18.7},
  {16, _, 18.4},
  {16.7, _, 18.7},
  {16.7, 20.2, 19.4},
  {17.7, 20.2, 19.9},
  {18.8, 21.1, 21.5},
  {20, 22.5, 24},
  {20.1, 23.8, 24.3},
  {21.1, 24.3, 25.6},
  {22.3, 24.9, 26.3},
  {22.9, 25.5, 26.2},
  {23.4, 25.5, 26},
  {22.2, 25.2, 26.2},
  {20.7, 23.9, 25},
  {19.8, 22.7, 24.8},
  {18.8, 21.4, 23},
  {18.7, 20.1, 20.2},
  {18.5, 19.8, 18.7},
  {16.8, 20.1, 17.9},
  {15.9, 19.5, 17.3},
  {15.5, 18.5, 16.7},
  {15.2, 18.4, 16.1},
  {16.1, 18.2, 16},
  {15.7, 17.4, 16},
  {15.7, 16.5, 15.5},
  {15.6, 16.5, 15.2},
  {18.3, 17.6, 16},
  {19.6, 18.9, 18.3},
  {19.6, 20.7, 21},
  {20.6, 21.8, 23.4},
  {22, 23.9, 25.4},
  {22.6, 25.4, 26.9},
  {22.7, 26.8, 27.4},
  {21.8, 24.6, 23.9},
  {21, 24.2, 25.4},
  {21.5, 22.3, 25.4},
  {20.8, 21.8, 25},
  {19.7, 20.9, 24.1},
  {19.7, 18.5, 23.6},
  {18.8, 17.8, 23},
  {18, 17.3, 21.2},
  {17.2, 17.1, 19.7},
  {15.5, 16.9, 17.9},
  {14.3, 16.1, 16.5},
  {14.4, 15.4, 15.9},
  {13.8, 14.8, 15.5},
  {13.3, 14.4, 15.2},
  {12.8, 14.1, 15.1},
  {12.3, 13.7, 14.7},
  {13.1, 13.7, 14.2},
  {14.3, 15, 14.7},
  {14.7, 15.5, 15.7},
  {14.6, 17.2, 17.3},
  {14.4, 17.6, 18.8},
  {14.7, 17.9, 18.8},
  {15, 17.5, 18.5},
  {16.2, 17.4, 18.4},
  {16.4, 17.5, 18.4},
  {16.4, 17.2, 18.9},
  {15.3, 17.5, 18.9},
  {14.1, 16.2, 19},
  {13.9, 15.8, 18.3},
  {13.9, 15.2, 17.4},
  {13.4, 15, 16.7},
  {13, 14.8, 16.5},
  {13.1, 14.7, 16.1},
  {13.1, 14.7, 15.8},
  {13.3, 14.8, 15.7},
  {13.4, 15, 15.7},
  {13, 14.8, 15.6},
  {12.5, 15, 15.3},
  {12.5, 14.7, 15.2},
  {12.2, 14.6, 15},
  {13, 14.6, 14.9},
  {14.1, 14.7, 15},
  {14.3, 15.2, 15.3},
  {16, 16.1, 16.5},
  {17.8, 18, 19.6},
  {19.3, 19.5, 22.2},
  {19.5, 20.3, 23.9},
  {20.2, 19.4, 25},
  {19.4, 22.1, 26.4},
  {19.9, 22.3, 25.3},
  {20.5, 21.8, 25.6},
  {18.8, 19.9, 24.2},
  {17.1, 18.8, 20.7},
  {16.6, 18.5, 19.4},
  {16.3, 17.7, 18.8},
  {15.8, 17, 18.4},
  {16, 16.8, 17.7},
  {16.2, 17, 17.3},
  {16.4, 17.1, 17.4},
  {15.9, 16.8, 17.1},
  {15.5, 16.7, 16.9},
  {15.2, 16.6, 16.7},
  {15.1, 16.3, 16.5},
  {14.8, 15.6, 16.3},
  {15.3, 16.1, 15.9},
  {16.3, 16.6, 15.9},
  {17.8, 17.7, 17},
  {18.4, 18.2, 18.1},
  {19.5, 18.7, 19.8},
  {20.6, 19.2, 21.7},
  {21.9, 20.7, 23.6},
  {22.1, 21.9, 25.7},
  {21.5, 23.1, 26.2},
  {22.1, 24.5, 24.4},
  {21.5, 24.8, 23.4},
  {20.7, 24.5, 23.7},
  {21.5, 24.4, 24.9},
  {18.6, 24.1, 24.9},
  {17.7, 21.5, 22.1},
  {16.6, 19.1, 19.8},
  {16.4, 18.5, 18.3},
  {16.9, 18.5, 17.4},
  {17.6, 18.5, 16.8},
  {17.2, 18.6, 16.7},
  {16.4, 18.4, 16.6},
  {15.9, 17.7, 16},
  {15.7, 17.2, 15.2},
  {15.6, 17, 14.7},
  {16.3, 16.4, 14.2},
  {18.1, 16.7, 14.5},
  {18.6, 18, 17},
  {19.3, 20.4, 20.5},
  {20.7, 22.7, 22.4},
  {22.4, 25.2, 24.9},
  {24.1, 26.7, 27.4},
  {25.2, 27.1, 28.6},
  {25.6, 28.5, 29.9},
  {25, 29, 29.2},
  {24.8, 28.5, 28.8},
  {24.3, 27, 28.2},
  {23.7, 25.5, 26.8},
  {22.1, 25, 26.8},
  {20.2, 24.2, 26.3},
  {19.3, 23.2, 23.5},
  {17.8, 22.6, 21.2},
  {17.1, 21.6, 20.2},
  {17.2, 20.6, 18.9},
  {17.7, 20.3, 18},
  {18.4, 20, 17.7},
  {18.5, 19.4, 17.9},
  {18.5, 18.8, 17.7},
  {17.8, 18.6, 17.5},
  {17.7, 18.5, 17.1},
  {21.1, 18.9, 17.5},
  {22.5, 20.2, 19.8},
  {22.9, 22, 22.3},
  {23.4, 23.6, 24.7},
  {24.1, 25.3, 26.6},
  {24.8, 26.7, 28.4},
  {25.3, 27.7, 28.9},
  {25.7, 28.3, 29.2},
  {25.6, 28.8, 28.7},
  {25.7, 29, 29},
  {25.6, 28.6, 29.3},
  {24.1, 27.8, 28.8},
  {22.9, 26.7, 27.9},
  {21.8, 24.8, 26.1},
  {19.7, 23.6, 22.4},
  {19.8, 22.5, 21},
  {19.9, 22.4, 20.3},
  {20, 22.4, 19.9},
  {19.3, 21.3, 19.3},
  {16.8, 19.8, 18.4},
  {15.9, 18.8, 18.1},
  {15.5, 17.9, 17.8},
  {15.5, 17.4, 17.1},
  {16.8, 17.9, 16.6},
  {19.8, 18.4, 17.1},
  {21.7, 19.4, 18.8},
  {21.6, 22.5, 21.2},
  {22.6, 25.3, 24.1},
  {24.1, 25.2, 26.7},
  {25.2, 26.5, 29},
  {25, 27.9, 31},
  {25.3, 27.6, 29.4},
  {25.1, 26.9, 28.8},
  {24.4, 26.8, 25.1},
  {20.1, 24.6, 19.9},
  {17.5, 22.8, 19.7},
  {18, 21.9, 19.7},
  {17.9, 20.6, 19.5},
  {17.4, 20.8, 19.1},
  {17.7, 19.3, 18.3},
  {16.7, 18.5, 17.2},
  {16.3, 17.7, 16.4},
  {15.5, 17.2, 16},
  {15.1, 16.5, 15.4},
  {15.2, 15.8, 15.1},
  {15.3, 15.4, 14.7},
  {14.1, 15.3, 14.6},
  {15.6, 15.4, 14.6},
  {18.3, 16, 14.5},
  {19.1, 17.3, 15},
  {19.4, 20.4, 16.4},
  {21.2, 20.8, 19.8},
  {22.3, 22.8, 23.7},
  {24.1, 24.9, 26.1},
  {24.3, 25.7, 27.7},
  {25.1, 27.2, 29.5},
  {24.5, 27.2, 29.5},
  {23.5, 26.8, 27},
  {22.2, 25.7, 22.1},
  {21.7, 25.5, 21},
  {20.8, 25, 20.8},
  {18.8, 22.5, 20.3},
  {17.7, 21.4, 18.6},
  {17.5, 21.1, 17.3},
  {17.6, 19.7, 16.7},
  {18.2, 18.7, 16.6},
  {18, 18.2, 16.5},
  {17.7, 17.6, 16.4},
  {18.4, 17.4, 16.4},
  {18.6, 17.4, 16.4},
  {16.7, 16.7, 15.8},
  {16.9, 16.4, 15},
  {19.9, 16.9, 15.2},
  {19.2, 18.6, 17},
  {20.3, 20.7, 20},
  {21.5, 23, 22.9},
  {22.7, 24.9, 25.2},
  {24.3, 25.3, 27.1},
  {25.2, 27.2, 28.9},
  {25.8, 28.5, 29.8},
  {25, 28.4, 29.1},
  {25.9, 28.3, 28.8},
  {24.8, 28.3, 27.8},
  {23.8, 27.1, 27.5},
  {22.4, 25.7, 26},
  {20.4, 18.9, 24.1},
  {19.8, 18, 21.4},
  {18.8, 17.3, 19.8},
  {18.5, 16.6, 19.2},
  {17.2, 16.4, 18.9},
  {17, 16.1, 18},
  {16.5, 16, 17.4},
  {16.3, 16.2, 16.4},
  {15.5, 15.7, 15.7},
  {15.6, 15.8, 15.1},
  {16.9, 15.9, 14.9},
  {18.5, 16, 15.4},
  {20.6, 17.2, 17.6},
  {21.3, 19.8, 20.7},
  {22.5, 22.1, 23.4},
  {23.3, 23.9, 25.7},
  {24.7, 26.1, 27.8},
  {24.9, 27.3, 28.2},
  {24.9, 28, 28.2},
  {24.8, 28.1, 28.4},
  {24.7, 28.1, 28.5},
  {24.6, 27.8, 28},
  {23.9, 26.7, 27.5},
  {22.6, 25.6, 26.8},
  {21.4, 24.2, 25.3},
  {20.7, 22.4, 22.7},
  {20.1, 22.3, 21},
  {19.5, 22, 20.3},
  {19.7, 21.3, 20.4},
  {19.7, 20.2, 20},
  {18, 19.8, 18.9},
  {19.1, 19.6, 18.4},
  {18.5, 20.6, 18.7},
  {18.4, 20.4, 18.9},
  {18.2, 20.2, 19},
  {18.3, 20.4, 19.5},
  {18, 20.8, 20.4},
  {17.8, 21.3, 21.7},
  {18.2, 22, 22.1},
  {20.1, 22.8, 24.1},
  {20.7, 23.6, 23.8},
  {21.2, 24.2, 24.6},
  {21.8, 24.8, 25.2},
  {21.7, 25.1, 25.5},
  {21.9, 25.2, 25.6},
  {21.8, 24.9, 25.4},
  {21.2, 24.3, 25.2},
  {19.4, 23.4, 24.6},
  {18.6, 21.4, 23.3},
  {17.7, 20.4, 20.9},
  {16.4, 19.4, 18.6},
  {16.5, 19.2, 18.4},
  {14.8, 19, 17.6},
  {14.3, 18.4, 16.4},
  {14.2, 17.8, 15.8},
  {13.8, 17, 15.3},
  {13.4, 16.9, 14.7},
  {13.3, 17.1, 14.4},
  {14.4, 17.3, 15},
  {15.8, 18.1, 16},
  {16.7, 18.9, 17.5},
  {17.9, 20.3, 20.9},
  {18.8, 21.4, 22.8},
  {20.4, 22.6, 23.9},
  {21, 23.8, 24.9},
  {22.5, 24.8, 25.8},
  {23.4, 25.6, 26.8},
  {24, 26.2, 27.3},
  {24.5, 26.5, 26.6},
  {23.9, 26, 26.3},
  {22.7, 25, 25.2},
  {20.7, 23.2, 24.2},
  {19.3, 21.9, 22.5},
  {17.6, 21, 19.4},
  {17.6, 20.3, 17.7},
  {15.3, 19.2, 16.7},
  {14.8, 19.1, 15.7},
  {14.3, 18.5, 14.7},
  {14.1, 17.3, 14.2},
  {13.6, 16.5, 13.6},
  {13.6, 15.7, 13.1},
  {13.4, 15.3, 12.7},
  {14.2, 15.3, 12.4},
  {17.9, 15.8, 13.1},
  {19.4, 16.7, 15.6},
  {19.8, 20.1, 19.4},
  {20.4, 21.8, 22.1},
  {21.8, 23.7, 24.8},
  {23, 25, 26.7},
  {24, 26.4, 27.5},
  {24.5, 27.3, 27.7},
  {24.7, 27.4, 27.7},
  {25.3, 27.5, 27.9},
  {25, 27.4, 27.5},
  {23.7, 26.4, 27.2},
  {20.8, 25, 26.6},
  {19.7, 23.2, 24.1},
  {17.2, 22, 19.8},
  {16.2, 21, 17.8},
  {15.8, 20.6, 16.7},
  {15.5, 19.7, 15.6},
  {15.2, 18.6, 14.9},
  {14.7, 17.8, 14.3},
  {14.2, 16.9, 13.7},
  {13.9, 16.3, 13.3},
  {14.2, 16, 12.8},
  {14.8, 16.6, 12.6},
  {19.3, 17, 13.1},
  {21.2, 18.5, 16.2},
  {21.6, 20.8, 20.2},
  {22.9, 22.3, 23},
  {24.8, 24.7, 25.9},
  {26.1, 27, 28.7},
  {27.3, 29.3, 30.9},
  {28, 30.2, 31.3},
  {28.1, 30.7, 30.7},
  {27.1, 30.3, 30.6},
  {26.4, 29.3, 30.1},
  {25.1, 28.3, 29.5},
  {24, 27.2, 29},
  {22.8, 25.8, 26.3},
  {19.4, 24.8, 21.7},
  {18.1, 23.4, 18.7},
  {17.5, 22, 17.4},
  {17.2, 20.9, 16.3},
  {16.8, 19.7, 15.5},
  {16.7, 19, 14.8},
  {16.2, 18.5, 14.2},
  {16.2, 18, 13.7},
  {16, 18.4, 13.1},
  {16.8, 18.5, 12.8},
  {21, 18.7, 13.2},
  {23, 20.5, 16.5},
  {23.6, 22.3, 21.2},
  {25.3, 23.8, 24},
  {26.9, 26.6, 27.2},
  {28.2, 29.1, 30.1},
  {29, 31, 32.3},
  {29.4, 31.7, 32.6},
  {29.2, 32.4, 32.7},
  {28.7, 32.2, 32.5},
  {28, 31.5, 31.6},
  {26.9, 30.6, 31.1},
  {25, 29.2, 29.9},
  {24.2, 27.3, 26.4},
  {21.3, 25.7, 21.4},
  {19.5, 24.9, 18.6},
  {18.8, 23.5, 17},
  {18.3, 22.1, 16.2},
  {18.1, 20.4, 15.7},
  {18.1, 20.1, 15.2},
  {17.8, 20.3, 14.5},
  {17.8, 20.1, 13.8},
  {17.2, 19.6, 13.5},
  {18.1, 19.3, 13.3},
  {22.1, 19.8, 14.1},
  {23.7, 21.3, 17.9},
  {24.6, 23.9, 22.1},
  {25.5, 24.7, 25.2},
  {27.5, 27.1, 28.7},
  {29, 29.6, 31.4},
  {29.9, 32.1, 34.1},
  {30.6, 33.1, 34.5},
  {30.2, 33.6, 34.4},
  {29.7, 33.3, 33.8},
  {28.8, 32.2, 33.2},
  {27.7, 31.1, 32},
  {25.7, 29.3, 30.4},
  {24.2, 27.9, 27.5},
  {22.5, 26, 22.2},
  {21, 25.1, 20.3},
  {20.9, 24, 19.1},
  {19.9, 22.6, 17.8},
  {19.4, 22.4, 16.9},
  {19.7, 22.2, 16},
  {19.5, 21.1, 16.3},
  {19.8, 20.4, 16},
  {18.5, 19.5, 15},
  {18, 19.4, 14.3},
  {20.8, 20.1, 14.9},
  {22.6, 21.3, 18.5},
  {23.3, 23.9, 22.3},
  {25.2, 26.5, 25.6},
  {27, 27.2, 28.5},
  {28.6, 29, 31.2},
  {29.1, 31, 32.8},
  {29.1, 32.2, 32.8},
  {28.6, 30, 32.9},
  {27.6, 29, 31.7},
  {26.2, 28.7, 27.6},
  {24.3, 27.8, 24.5},
  {23.8, 26, 24},
  {22.3, 24.8, 22.1},
  {21.6, 23.4, 21.5},
  {21.7, 23.4, 20},
  {21.6, 22.1, 19.1},
  {20.5, 20.3, 18.2},
  {19.2, 19.4, 17.5},
  {18.5, 19.1, 16.7},
  {17.6, 18.4, 16.2},
  {16.8, 18.1, 15.6},
  {17.6, 17.9, 14.8},
  {17.5, 17.8, 14.8},
  {20.2, 18.1, 15.3},
  {21.4, 19.2, 17.8},
  {22.2, 20.8, 21.4},
  {24, 23.4, 24.9},
  {25.3, 25.5, 28},
  {27.3, 27.3, 30.5},
  {28.8, 28.6, 32.5},
  {29.7, 29.6, 32.7},
  {26.7, 29.2, 28.5},
  {25.4, 28.9, 26.9},
  {24.8, 28.2, 26.1},
  {24.7, 25.3, 25.6},
  {23.7, 23.9, 24.9},
  {21.4, 22.5, 23},
  {20.3, 22.1, 20.4},
  {21.6, 22.5, 18.9},
  {21.2, 22.7, 18.9},
  {21.4, 22.1, 19.2},
  {20.5, 21.2, 19.1},
  {20.5, 21.1, 18.8},
  {19.3, 20.5, 18.7},
  {17.9, 19.2, 18.4},
  {17.8, 19, 16.8},
  {17.7, 18.8, 16.4},
  {19.9, 18.7, 16.4},
  {21, 19.5, 19.3},
  {22.3, 22.3, 23.6},
  {23.6, 25, 26.2},
  {25, 25.9, 28.3},
  {26.9, 27.6, 30.8},
  {28, 29.2, 32.6},
  {28.4, 30.9, 32.6},
  {28.1, 31.6, 32.6},
  {27.7, 31.3, 32.1},
  {27, 30.4, 31},
  {26, 29, 30.4},
  {24.6, 27.7, 29.7},
  {22.8, 26.2, 28},
  {22.5, 24.8, 24.6},
  {22.6, 24.1, 22.5},
  {21.6, 24.1, 22},
  {20.9, 23.8, 21.7},
  {20.4, 21.3, 18.3},
  {20.4, 20.7, 17.7},
  {19.3, 19.5, 17.6},
  {18.1, 18.3, 17.3},
  {17.6, 18.2, 16.8},
  {17.5, 17.9, 16.5},
  {21, 18.2, 16.6},
  {21.1, 19.5, 17.7},
  {21.8, 22.2, 19.7},
  {23.7, 23, 22.3},
  {25.5, 25.2, 25.4},
  {26.5, 27.8, 27.6},
  {27.7, 29.3, 29.7},
  {28.2, 30.8, 31.4},
  {27.9, 31.4, 31.6},
  {28.1, 30.8, 30.5},
  {25.8, 30.2, 28.7},
  {24.7, 28.5, 26.8},
  {23.7, 27.4, 24.9},
  {22.8, 25.7, 22.8},
  {20.8, 24.8, 21.3},
  {20.4, 24.4, 20.4},
  {20.9, 24.3, 19.8},
  {20.7, 21.9, 18.9},
  {20.8, 17.6, 18.4},
  {21, 17.4, 18.4},
  {17.9, 17.1, 18.8},
  {16, 16.8, 18.8},
  {15.8, 16.5, 18.4},
  {16.2, 16.3, 17.8},
  {18, 16.5, 17.9},
  {19.3, 16.9, 19.2},
  {20.3, 18.6, 21.7},
  {21.9, 20.8, 24.1},
  {23.8, 22.9, 26.2},
  {25.3, 24.8, 28.4},
  {26.8, 27.4, 30.1},
  {27.6, 29.7, 32.1},
  {27.1, 30.2, 31.9},
  {23.8, 28, 29.1},
  {22.2, 25.3, 27.5},
  {22.6, 24.8, 26},
  {22.2, 23.5, 25.3},
  {21.1, 21.3, 23.7},
  {20.8, 20.7, 22.5},
  {20.7, 22.1, 21},
  {20.7, 20.9, 20.4},
  {20.6, 19.2, 20.3},
  {19.2, 19.4, 19.9},
  {18.7, 19.2, 19.5},
  {18.2, 18.9, 18.7},
  {17.9, 18.6, 18.6},
  {17.3, 18.3, 18.2},
  {17, 18.4, 17.7},
  {19.1, 18.5, 17.4},
  {20.2, 19.2, 19},
  {21.4, 21.1, 21.1},
  {22.9, 23.8, 24.2},
  {24.5, 24.7, 26.7},
  {26.6, 26.2, 28.9},
  {27.5, 28.6, 30.7},
  {28.3, 30, 32},
  {28.3, 30.8, 31.9},
  {28.1, 29.9, 32.3},
  {27.5, 30.1, 31.1},
  {25.9, 28.7, 31.1},
  {24.1, 26.8, 29.2},
  {22.1, 25.4, 26.3},
  {20.7, 23.9, 23.2},
  {20.1, 23.7, 21.8},
  {19.2, 22.8, 21},
  {19, 19.4, 19.9},
  {19.8, 18, 19.5},
  {19.4, 16.8, 21.9},
  {17.6, 16.5, 22.2},
  {15.8, 16.8, 20.3},
  {15.1, 16.5, 18.1},
  {14.7, 16.8, 16.8},
  {18.5, 17, 16.7},
  {20.3, 17.5, 18.7},
  {20.4, 19.3, 21.9},
  {21.3, 21.6, 24.4},
  {23.4, 23.4, 26},
  {25.3, 24.6, 28.2},
  {26.5, 26.6, 29.7},
  {27.3, 28.3, 30.2},
  {28, 26.9, 27.9},
  {26.2, 26.6, 20.6},
  {24.1, 25.4, 18.2},
  {21.3, 23.5, 18},
  {17.9, 19, 17.7},
  {18.8, 16.6, 17.5},
  {17, 16, 17.5},
  {17.5, 15.9, 16.8},
  {17.4, 15.8, 16.4},
  {17.1, 15.8, 16.4},
  {17.2, 16, 16.2},
  {15.8, 15.8, 15.8},
  {15.5, 16, 15.4},
  {15.2, 16.1, 15.2},
  {14.8, 16.1, 15.2},
  {15.3, 16.4, 15.2},
  {16.1, 16.4, 15.4},
  {16.3, 16.4, 15.7},
  {16.9, 16.3, 16.1},
  {17.9, 16.6, 17.4},
  {18.5, 16.7, 20},
  {18.8, 17.4, 21.8},
  {20, 18.2, 22.6},
  {20.9, 19.3, 23.2},
  {21.4, 20.1, 25.1},
  {22.2, 20.4, 25.9},
  {21.4, 21.7, 26.3},
  {20.3, 22.6, 24.9},
  {20.2, 21, 25.4},
  {18.8, 20.2, 22.3},
  {16.9, 19.5, 19.6},
  {16.5, 18.6, 18.5},
  {15.6, 18.4, 17.4},
  {15.5, 17.6, 16.5},
  {14.7, 17.1, 15.7},
  {14.7, 16.7, 15.2},
  {15.5, 16.4, 14.6},
  {14.6, 16.4, 14.1},
  {14.9, 16.2, 13.8},
  {15.1, 16, 13.6},
  {18, 16.5, 14},
  {19.4, 17.9, 15.3},
  {20.7, 20, 17},
  {22.1, 23, 21},
  {23.7, 25.6, 24.2},
  {25.6, 27.4, 27.2},
  {26.4, 27.2, 29.4},
  {26.4, 28.9, 30.1},
  {25.6, 29.5, 29.3},
  {26.2, 29.1, 29.1},
  {26, 28.5, 28.9},
  {24.6, 27.2, 28.3},
  {23.3, 25.8, 27.3},
  {22.8, 24.3, 26},
  {21.9, 23.4, 22.5},
  {21.2, 23, 20.7},
  {20.2, 22.1, 19.4},
  {19.3, 21.1, 19},
  {19, 20.8, 18.3},
  {18.5, 20.3, 17.9},
  {18.2, 19.4, 17.6},
  {19.2, 17.9, 17.6},
  {18.3, 17.9, 17.8},
  {17.2, 18.2, 18.3},
  {17.6, 18.2, 18.3},
  {19.6, 18.5, 19.4},
  {20.7, 20.8, 21.8},
  {21.9, 22.9, 24.6},
  {23.1, 24.3, 26.4},
  {25.2, 25.1, 28.2},
  {26.5, 26.9, 29},
  {27.6, 26.6, 30.8},
  {27.5, 28.5, 29},
  {20.2, 28.3, 21},
  {19.2, 26.6, 21},
  {19.8, 26.4, 20.9},
  {19.7, 24.9, 20.3},
  {19.3, 21.9, 20},
  {18.8, 18.6, 19.4},
  {18.3, 18.3, 18.7},
  {18.9, 17.9, 18.2},
  {18.9, 18, 17.9},
  {18.2, 17.8, 17.8},
  {17.3, 17.2, 17.8},
  {16.4, 16.8, 17.8},
  {16, 16.7, 17.5},
  {15.4, 16.1, 17.1},
  {15.2, 15.8, 17.1},
  {16.3, 16.5, 17.1},
  {16.3, 16.8, 17.1},
  {16.3, 16.8, 17.3},
  {15.8, 16.7, 17.2},
  {16.1, 17.5, 17.7},
  {17, 18.3, 18.3},
  {19.7, 19.9, 20.8},
  {21.7, 21.7, 23.8},
  {22.4, 21.3, 26.1},
  {22.3, 19.5, 25.3},
  {21.4, 18.9, 22.8},
  {19.4, 18.6, 21.2},
  {18.6, 18, 21.4},
  {18, 17, 20.8},
  {17.3, 16.1, 19.7},
  {16.9, 16.6, 18.8},
  {16.6, 16.8, 18.6},
  {16.3, 16.8, 18.1},
  {15.4, 16.7, 17.5},
  {15, 16.9, 16.7},
  {15, 16.9, 16.2},
  {14.8, 16.6, 15.6},
  {14.5, 16.1, 15.3},
  {14.1, 15.9, 15.2},
  {15.9, 15.5, 15.6},
  {17.5, 15.4, 16.5},
  {17.9, 16.9, 18},
  {18.3, 18.6, 19.9},
  {19.7, 21.3, 22.4},
  {20.9, 23.1, 24.7},
  {20.8, 22.9, 26.2},
  {21.9, 23.6, 25.4},
  {21.7, 23.9, 24.2},
  {18.8, 23.4, 23.1},
  {17.8, 22.1, 22.2},
  {17.3, 21.3, 22.3},
  {16.5, 20, 22.1},
  {16.1, 18.9, 21.1},
  {15.4, 18.4, 19.6},
  {15.3, 18.2, 19.1},
  {15.3, 17.9, 18.5},
  {15.4, 17.8, 18.2},
  {15.2, 15.7, 18.2},
  {14.9, 14.2, 18},
  {14.5, 13.9, 17.7},
  {12.7, 13.9, 17.3},
  {12.3, 13.5, 16.2},
  {12.2, 13.2, 15.6},
  {12.2, 13.5, 15.4},
  {12.4, 13.5, 15.1},
  {12.6, 13.8, 15.1},
  {12.8, 13.6, 15.3},
  {13, 13.7, 15.2},
  {12.7, 13.4, 15.1},
  {12.5, 12.4, 15},
  {12.7, 11.4, 14.7},
  {12.3, 12.7, 15.8},
  {12.9, 14.7, 17.8},
  {14.2, 15.8, 19.2},
  {14, 15.9, 19.1},
  {13.8, 14.9, 17.5},
  {12.1, 14, 16.6},
  {12, 14.1, 14.6},
  {12.3, 13.9, 13.9},
  {12.9, 14.9, 10.4},
  {11.8, 15.3, 10.4},
  {10.9, 14.3, 10.3},
  {10.2, 14, 10.1},
  {10.2, 14.6, 9.9},
  {9.9, 15.7, 9.8},
  {9.8, 14.8, 9.8},
  {10.5, 14, 9.1},
  {11.4, 13.1, 9},
  {12.9, 14.9, 9.1},
  {13.7, 15.4, 9.5},
  {14.2, 15.7, 11},
  {14.5, 16.5, 10.9},
  {15.2, 17.2, 12.4},
  {15.8, 16.5, 13.9},
  {16.9, 17.8, 15.4},
  {17.5, 20.4, 16.5},
  {18.1, 20.9, 17.3},
  {18.1, 21.1, 18.2},
  {15, 20.3, 17},
  {15.3, 17.9, 14.4},
  {13.1, 14.9, 12.1},
  {11.9, 13.4, 10.8},
  {11.5, 12.8, 9.5},
  {10.7, 13.1, 8.9},
  {10.5, 13.3, 8.3},
  {10.1, 12.8, 8.2},
  {9.9, 11.9, 8.4},
  {9.3, 10.8, 7.6},
  {9.2, 10.4, 6.9},
  {9.3, 9.7, 6.8},
  {9, 9.6, 7.1},
  {10.4, 11.8, 7.6},
  {13.6, 14.1, 11.4},
  {15.6, 15.5, 15},
  {16.4, 15.8, 16.3},
  {17.3, 18.3, 17},
  {19.1, 19.8, 18},
  {19.3, 20.2, 18.9},
  {20.2, 22.7, 19.5},
  {20.3, 23.7, 20.6},
  {19.3, 23.8, 20.6},
  {18.9, 23.7, 20.7},
  {17.7, 22.4, 20.2},
  {17.2, 18.9, 15.8},
  {16.2, 15.8, 14.6},
  {15.4, 14.4, 13.1},
  {14.4, 13.4, 11.5},
  {12.6, 13.1, 10.7},
  {12.6, 12.8, 10},
  {12.2, 12.8, 9.2},
  {11.7, 13.1, 8.9},
  {11.2, 12.7, 8.4},
  {10.9, 12, 9.2},
  {10.8, 12.1, 10},
  {11.3, 12.5, 10.2},
  {13.8, 13.4, 10.8},
  {14.6, 15.2, 12},
  {17, 18.5, 15.4},
  {18, 19.9, 17.2},
  {18.9, 21.6, 19.5},
  {20.5, 22.7, 20},
  {21.5, 23.7, 21},
  {21.2, 24.7, 20.7},
  {15.5, 23.4, 21.2},
  {14.3, 23.2, 20.9},
  {15.6, 22, 21.1},
  {17.9, 20.8, 20},
  {14.4, 19.4, 18.4},
  {13.5, 16.1, 15.7},
  {13.5, 15.5, 14.3},
  {13.7, 15.7, 12.8},
  {13.5, 15.4, 11.8},
  {12.6, 15.3, 11.3},
  {12.7, 15.2, 10.9},
  {13.1, 15.8, 10.7},
  {13.4, 15.8, 10.5},
  {13.2, 15.1, 10.9},
  {13.5, 15.3, 11},
  {13.1, 15.1, 10.6},
  {14, 15.1, 10.9},
  {14.9, 16.4, 15.2},
  {16.1, 19, 18.1},
  {17.9, 21, 19.1},
  {19.8, 21.5, 19.7},
  {20.5, 21.1, 20},
  {20.6, 23.1, 20.4},
  {21.2, 23.7, 20.6},
  {22, 23.6, 20.8},
  {22.2, 23.8, 20.7},
  {22.1, 23.6, 20.9},
  {20.5, 23.2, 19.5},
  {17.3, 22, 18.7},
  {16.6, 20.8, 14.9},
  {15.9, 18.2, 13.2},
  {15.5, 16.3, 12.8},
  {15.5, 15.5, 11.4},
  {14.9, 16.1, 11},
  {14.7, 16.2, 10.2},
  {14.1, 16.4, 9.9},
  {13.5, 15.9, 9.3},
  {12.3, 14.7, 9.1},
  {12.2, 14.8, 8.9},
  {11.7, 15.9, 8.7},
  {15.5, 16, 9.4},
  {18.1, 16.9, 13.2},
  {18.6, 17.8, 15.1},
  {19.5, 20.1, 16.3},
  {20.9, 22.7, 17},
  {20.9, 22.4, 18.2},
  {21.5, 22.8, 19},
  {22, 22.9, 20.8},
  {21.7, 23.7, 21.6},
  {22.2, 24.7, 22},
  {22.5, 24.3, 21.5},
  {21.3, 23.7, 20.7},
  {18.1, 22.4, 16.1},
  {17.9, 20.5, 14.3},
  {18, 18.3, 13},
  {16.4, 17.5, 11.9},
  {15.3, 18, 11.6},
  {15.5, 15.4, 10.8},
  {15.4, 14.9, 10.8},
  {13.9, 14.2, 10.8},
  {14.1, 13.2, 10.7},
  {13.9, 13.7, 9.6},
  {12.6, 13.2, 8.7},
  {12.4, 13.5, 8.5},
  {14, 14.4, 9.2},
  {16.3, 15.6, 12.1},
  {16.5, 16.6, 15.1},
  {18.5, 19.2, 18.6},
  {18.9, 21.6, 19.6},
  {19.8, 22.3, 17.2},
  {20.4, 22.2, 18.9},
  {20, 20.9, 19.3},
  {19.7, 19.5, 20.8},
  {18.9, 17.3, 19.1},
  {17.3, 14.5, 16.5},
  {15.2, 13.5, 14.5},
  {13.4, 13.1, 13.7},
  {12.3, 12.5, 12.9},
  {11.9, 11.7, 12.1},
  {11.7, 11.5, 11.6},
  {11.8, 11.9, 11.3},
  {11.7, 12, 11.4},
  {11.5, 11.8, 11},
  {11.3, 11.1, 11},
  {11.2, 11, 10.9},
  {10.9, 10.8, 10.3},
  {10.8, 10.7, 10.7},
  {10.4, 10.6, 10.7},
  {11.4, 11.4, 10.6},
  {13.8, 12.6, 12.5},
  {14.6, 14.8, 14.6},
  {14.8, 16.2, 16},
  {17.4, 18.1, 18.5},
  {18.4, 20.3, 19.8},
  {18.6, 20.8, 19.9},
  {16.6, 20.4, 18.6},
  {18.6, 21.9, 19},
  {18.4, 19.5, 20.1},
  {18.3, 18, 18.9},
  {17.8, 15.8, 17.6},
  {16.6, 14.7, 14.6},
  {13.1, 14, 13.4},
  {13.2, 13.7, 12.3},
  {12.7, 13.3, 11.6},
  {11, 12.7, 11},
  {10.9, 12.8, 10.2},
  {10.7, 12.6, 9.1},
  {10.7, 11.9, 8.6},
  {10.5, 11.7, 8.3},
  {10.3, 11.2, 8.3},
  {10.3, 10.9, 8.4},
  {10.3, 11, 8.6},
  {10.7, 11.2, 9.1},
  {12.1, 12.3, 10.5},
  {13, 13.5, 12.6},
  {14.6, 15.3, 14.3},
  {15.8, 15.7, 15.4},
  {15.7, 16.8, 15.6},
  {14.8, 17.4, 18.2},
  {14.4, 16.8, 16.9},
  {15.4, 17.9, 11.1},
  {15.2, 17.4, 10.4},
  {15.4, 15.7, 11.1},
  {14.7, 13, 11.9},
  {13.4, 12.1, 11.6},
  {12.2, 11.8, 10.7},
  {11.4, 11.7, 10.5},
  {10.6, 11.3, 10.4},
  {10, 11.2, 10},
  {9.7, 11.1, 9.8},
  {9.6, 10.9, 9.1},
  {9.6, 10.5, 8.9},
  {9.5, 10.3, 8.8},
  {9.5, 10.3, 8.7},
  {9.2, 10.4, 8.7},
  {8.9, 10.5, 8.8},
  {9.4, 11, 9.2},
  {9.9, 11.2, 9.5},
  {11, 11.9, 10.7},
  {12.4, 13.9, 12.6},
  {13.8, 15.7, 15},
  {14.8, 16.9, 15.6},
  {12.8, 17.6, 14},
  {12.6, 14.7, 11.6},
  {12.3, 12.7, 10.9},
  {11.6, 13.3, 10.2},
  {10.6, 12.1, 9.4},
  {9.9, 11.9, 9.4},
  {9.5, 12.5, 9.2},
  {8, 10.6, 8.8},
  {6.9, 8.3, 8},
  {6.6, 7.5, 7.5},
  {6.3, 7.2, 6.7},
  {6.2, 7.3, 5.7},
  {6, 7.4, 5.2},
  {5.7, 7.2, 4.8},
  {6, 6.8, 4.6},
  {5.8, 6.3, 4.4},
  {6, 5.8, 4.3},
  {6.9, 6.6, 4.1},
  {7.9, 8.2, 5.3},
  {9.6, 9.5, 7.4},
  {11, 11.4, 10.9},
  {12.1, 13, 13.5},
  {13, 14.8, 15.1},
  {14.8, 16.4, 16.4},
  {15.4, 17.7, 17.1},
  {14.3, 18, 17.1},
  {13.2, 17.9, 16.7},
  {12, 17.9, 14.6},
  {12.5, 17.7, 15},
  {13.5, 16.6, 14.9},
  {12.9, 15.9, 12.5},
  {12.1, 12.4, 11.6},
  {11.5, 11.8, 10.7},
  {11.2, 11.3, 9.8},
  {11.2, 11.2, 9.3},
  {11.5, 11.7, 9.7},
  {10.5, 11.9, 9.8},
  {9.3, 11.8, 9.5},
  {8.9, 10.8, 9.3},
  {8.2, 10.7, 9.1},
  {8.8, 10.7, 8.9},
  {8.8, 10.7, 8.7},
  {9.1, 10.6, 8.9},
  {9.7, 11.1, 9.2},
  {10.3, 11.3, 9.5},
  {12.2, 12, 10.3},
  {14, 13.3, 11.2},
  {15.2, 15.1, 13.1},
  {16.1, 16.5, 14.6},
  {16.2, 18, 16.4},
  {14.9, 14.9, 14.8},
  {15.1, 13.7, 17.4},
  {15.4, 14.5, 17.4},
  {13.5, 13.8, 15.3},
  {11.1, 13.6, 13.2},
  {9.9, 11.8, 12.2},
  {10.9, 10.4, 11.5},
  {11.8, 10.7, 9.8},
  {10.9, 10.4, 8.8},
  {10.1, 9.4, 7.8},
  {9.4, 8.8, 7.2},
  {9, 8.6, 6.8},
  {8.6, 8.9, 6.4},
  {8.5, 8.3, 6.1},
  {8.1, 8.5, 5.8},
  {8.1, 8.8, 5.7},
  {9.4, 9.9, 5.9},
  {10.9, 11.2, 7.7},
  {12.6, 13.3, 12.2},
  {14.6, 15.5, 15.5},
  {16.2, 17.1, 16.6},
  {17.2, 18.2, 17.9},
  {18.2, 19.6, 19.2},
  {18.6, 20.7, 19.8},
  {18.8, 20.8, 21},
  {18.4, 20.5, 21.1},
  {17.4, 19.5, 20},
  {16.2, 19, 17.4},
  {15.3, 17.8, 15.2},
  {14.2, 16.2, 13.8},
  {12.4, 15.2, 12.5},
  {11.6, 13.4, 10.9},
  {12, 13.7, 10.2},
  {12.2, 14.2, 10.1},
  {12.5, 14.3, 10.7},
  {13.3, 14.4, 11},
  {12.6, 13.8, 10.9},
  {12.2, 13, 10.6},
  {12.1, 12.7, 10.6},
  {12, 12.6, 10.6},
  {12, 12.5, 10.7},
  {12.4, 12.9, 10.6},
  {12.1, 13.3, 11.6},
  {12, 13, 11.7},
  {12, 13.2, 11.7},
  {12.7, 13.6, 12.6},
  {13.5, 14.8, 13.1},
  {13.5, 15.1, 14.5},
  {14.5, 15, 15.2},
  {14.3, 15.4, 16.5},
  {13.7, 15, 15.7},
  {13.6, 14.7, 14.3},
  {13.4, 14.4, 13.9},
  {13.2, 14.2, 13.3},
  {13.3, 14, 12.9},
  {13.3, 13.9, 12.6},
  {13.5, 13.9, 12.3},
  {13.7, 13.8, 12.3},
  {13.5, 13.8, 12.6},
  {13.2, 13.6, 12.2},
  {13.4, 13.6, 12},
  {13, 13.2, 12.1},
  {13.1, 12.7, 11.8},
  {13.7, 12.9, 12},
  {14, 13.5, 12.3},
  {15.8, 14.3, 13},
  {17, 15.9, 15.4},
  {18.6, 17.5, 18},
  {19.2, 19.2, 18.9},
  {19.6, 19.9, 20.9},
  {20.4, 21.1, 21.9},
  {20, 21.7, 21.1},
  {20.4, 21.9, 19.8},
  {20.9, 21.9, 21.6},
  {21.4, 21.3, 20.9},
  {19.8, 20.9, 20},
  {18.7, 20, 17.7},
  {17.4, 19.4, 16.6},
  {16.1, 17.7, 15.9},
  {15.4, 18.1, 14.9},
  {16.5, 18.3, 14.7},
  {16.4, 17.6, 14.7},
  {17.3, 18, 14.5},
  {17.1, 18.3, 14.3},
  {16.5, 17.6, 14.1},
  {16.1, 16.6, 13.6},
  {15.6, 15.8, 13.5},
  {15.5, 15.8, 13.5},
  {15.6, 16, 13.6},
  {16, 17.5, 14.3},
  {16.7, 18.2, 15.1},
  {17.8, 18.2, 16.2},
  {19.7, 21.9, 19.7},
  {20.9, 24, 21.5},
  {21.7, 24.6, 22.8},
  {21.7, 25.3, 23.9},
  {21.5, 24.8, 22.8},
  {21.7, 25.2, 22.9},
  {21.5, 24.8, 23.4},
  {20.7, 22.7, 21.7},
  {18.3, 19.3, 17.1},
  {16.7, 15.7, 15},
  {15.2, 15, 14},
  {15.3, 14.4, 13.4},
  {15.2, 14.1, 12.9},
  {15.5, 14.4, 12.5},
  {16, 15.2, 12.6},
  {16, 15.4, 12.7},
  {15.6, 14.6, 13.2},
  {15.2, 14.4, 13.7},
  {15.7, 14.3, 13.3},
  {15, 14.3, 12.9},
  {14.8, 14.8, 13.6},
  {16.6, 16, 14.4},
  {16.5, 18.3, 17.1},
  {16.6, 18.8, 19.5},
  {16.8, 18.1, 19.5},
  {19, 20.2, 21.4},
  {19.2, 21.6, 22.4},
  {18.5, 22, 21.7},
  {16.9, 19.9, 18.6},
  {19.2, 20.5, 17.6},
  {20.7, 21.8, 17.5},
  {18.6, 20.1, 17.8},
  {16.9, 18.6, 17.5},
  {15.9, 17.2, 15.9},
  {15.9, 16.3, 15.3},
  {15.6, 15.7, 15.4},
  {14.8, 15.2, 14.9},
  {14.5, 14.8, 14.2},
  {14.5, 14.4, 13},
  {13.8, 14.1, 12.1},
  {13.8, 13.8, 11.9},
  {13.6, 13.5, 11.6},
  {13.4, 13.2, 11.3},
  {13.3, 13.2, 10.7},
  {14, 14.4, 11.4},
  {16.8, 16.1, 13},
  {18.2, 18.7, 16.3},
  {19.4, 20, 20.3},
  {20.5, 21, 21.6},
  {20.9, 22, 22.7},
  {21.3, 23.2, 23.7},
  {21.5, 24.2, 23.7},
  {21.4, 25, 23.9},
  {20.6, 24.1, 20.6},
  {18, 18.3, 14.2},
  {18.6, 17.3, 14.8},
  {17.3, 16, 13.3},
  {15.3, 14.4, 12.3},
  {14.4, 13.2, 11.8},
  {13.7, 12.4, 11.2},
  {12.7, 11.9, 10.7},
  {11.7, 11.4, 10.3},
  {12.1, 11.1, 9.5},
  {11.9, 11, 9.3},
  {11.4, 10.7, 9.1},
  {11.6, 10.6, 8.9},
  {12.3, 10.6, 8.1},
  {12.3, 11.3, 8},
  {12.3, 12, 9.1},
  {13.2, 13, 10.1},
  {14.8, 15.1, 12.9},
  {16.6, 17.4, 16.8},
  {17.4, 19.3, 18.9},
  {18.9, 21, 20.5},
  {20.3, 22, 21},
  {20.1, 22.2, 21.4},
  {18.2, 22.2, 20.5},
  {19.4, 22.8, 21.3},
  {19.3, 22.9, 21.7},
  {18.2, 21.5, 20.5},
  {16.9, 17.8, 16.7},
  {16.3, 14.8, 14.3},
  {15.6, 13.8, 12.8},
  {14.6, 13.3, 12},
  {13.5, 13, 11.7},
  {13.4, 12.7, 11.3},
  {14.1, 13.3, 10.5},
  {14.5, 14, 10.4},
  {14.3, 14.2, 10.7},
  {13.6, 13.7, 10.7},
  {13.1, 12.6, 10.2},
  {13.7, 12.9, 10.1},
  {14.4, 14, 10.1},
  {15.6, 16, 11.9},
  {16.1, 17.7, 15.8},
  {17.2, 18.5, 18.6},
  {19.1, 20.2, 19.8},
  {19.4, 21.3, 19.6},
  {20.4, 22.4, 20.1},
  {20.5, 23.1, 22.3},
  {20.7, 22.1, 22.9},
  {20.8, 20.9, 23.2},
  {20, 22.5, 20.9},
  {18.7, 20.6, 20.9},
  {17.4, 17.8, 18.1},
  {15.5, 15.7, 15.2},
  {14.9, 15, 13.9},
  {14.5, 14.7, 13.2},
  {15.5, 15.2, 13.4},
  {15.7, 14.8, 13},
  {15.7, 14.8, 12.4},
  {16, 14.9, 12.2},
  {15.7, 15, 12},
  {15.1, 15, 11.7},
  {14.4, 14.7, 11.9},
  {14.1, 14.5, 12},
  {14.6, 14.7, 12.4},
  {15.9, 16.5, 13.6},
  {16.9, 17.6, 16.4},
  {18.1, 18.6, 18.5},
  {18.9, 20, 20},
  {19.7, 21.4, 21.2},
  {20.5, 22.1, 21.9},
  {19.9, 22.9, 22.9},
  {19.8, 22.8, 23.3},
  {20, 22.5, 23.3},
  {19.2, 21.5, 22.6},
  {19, 20.7, 20.8},
  {18.2, 19, 19.3},
  {17.6, 17.6, 17.9},
  {16.2, 17, 16.5},
  {15.7, 16.1, 15.8},
  {16.1, 16.5, 14.5},
  {16.6, 18.1, 14},
  {16.2, 17.2, 13.7},
  {15.8, 16.2, 13.5},
  {15.7, 16, 12.7},
  {14.3, 15.6, 12.4},
  {14.1, 15, 12.1},
  {14.5, 14.3, 12.1},
  {15.3, 15.1, 12.8},
  {16.1, 16.7, 14.8},
  {16.3, 17.6, 16.3},
  {15.9, 18.6, 18.5},
  {16.7, 19.4, 19.1},
  {17.9, 21.1, 21.3},
  {19.7, 22.4, 21},
  {20, 23.2, 21.2},
  {19.6, 22.1, 22.1},
  {19.2, 21.2, 20.9},
  {18.2, 20.8, 20.2},
  {17.1, 19.7, 19},
  {16.6, 17, 17.8},
  {15.7, 14.5, 16.9},
  {15, 14.4, 15.3},
  {14.7, 14.5, 14.2},
  {13.6, 14.9, 14.1},
  {12.7, 14.1, 14.1},
  {12.4, 14, 13.6},
  {12.5, 13.2, 12.5},
  {12.5, 12.8, 11.8},
  {11.8, 12.3, 11.5},
  {10.2, 11.3, 11.1},
  {9.4, 10.4, 11.1},
  {9.6, 10.8, 10.7},
  {11.4, 14.2, 11.9},
  {13.3, 16, 15.6},
  {14.8, 16.8, 17.1},
  {16, 17.8, 18.8},
  {17.1, 17.7, 20.1},
  {18.5, 18.6, 19.8},
  {18.9, 20.9, 21.3},
  {19.1, 18.8, 21.5},
  {18.5, 18.8, 20.6},
  {16.6, 18.3, 18.6},
  {14.4, 17.6, 17.8},
  {13.2, 16.1, 15.6},
  {12.9, 14.3, 13.2},
  {12.5, 13.6, 13},
  {12.5, 12.6, 12.3},
  {12.8, 13, 11.5},
  {13.3, 11.9, 11.8},
  {12.6, 13.1, 11.2},
  {12.2, 12.4, 10.8},
  {12, 11.9, 10.6},
  {11.3, 11.9, 10},
  {10.3, 11.6, 9.7},
  {10.2, 11.2, 9.5},
  {10.4, 11.1, 9.7},
  {12.3, 13.3, 10.9},
  {13, 15.4, 13.6},
  {16.2, 17.1, 15.8},
  {17.2, 18.6, 18},
  {18, 19.7, 19.5},
  {18.6, 19, 20.3},
  {18.3, 21.5, 21.2},
  {17.2, 20.9, 21.3},
  {17.7, 20.4, 21.2},
  {17.7, 19.7, 19.8},
  {17.1, 19.2, 18.7},
  {16.2, 17.4, 17.1},
  {14.9, 16.8, 15.5},
  {13.7, 15.3, 14},
  {14.4, 16.6, 13.8},
  {14.7, 16.1, 13.4},
  {14.6, 15.8, 13.1},
  {13.9, 12.5, 9.1},
  {11.2, 10.4, 9.2},
  {10.3, 10.4, 9.3},
  {9.8, 10.2, 8.9},
  {9.3, 9.9, 8.7},
  {8.6, 8.9, 8.1},
  {8.7, 9.1, 8.3},
  {11.1, 10.7, 9.1},
  {12.9, 13, 12.2},
  {14.2, 15.1, 15.1},
  {15.3, 16.9, 16.7},
  {16.8, 18.1, 18.6},
  {17.6, 19.6, 19},
  {18.6, 20.7, 19.6},
  {19.2, 21.5, 20.8},
  {18.6, 20.5, 20.7},
  {17.2, 17.6, 18.3},
  {16.4, 17.5, 16.6},
  {14.8, 14.4, 13.7},
  {13.2, 12.7, 12.6},
  {13, 12.4, 12},
  {12.6, 11.8, 11.2},
  {12.2, 11.5, 10.4},
  {11.7, 11.1, 9.7},
  {11.3, 10.5, 9.3},
  {10.9, 10.2, 8.7},
  {10.9, 9.6, 8.4},
  {10.5, 9.2, 7.6},
  {10.1, 8.9, 7.4},
  {9.7, 8.8, 7.1},
  {10.9, 10.6, 7.9},
  {13.1, 12.6, 9.8},
  {14.4, 13.3, 11.5},
  {14.3, 14.7, 13.3},
  {14.8, 14.6, 14.1},
  {15.9, 14.9, 14.4},
  {15.8, 15.7, 15.6},
  {16.6, 17, 17.3},
  {16.4, 18, 16.8},
  {15.7, 17.7, 16.4},
  {16.5, 17, 15},
  {16.5, 17.5, 13.8},
  {15.8, 17.5, 13},
  {15.2, 16.8, 12.4},
  {15, 15.6, 12.3},
  {15.2, 15.5, 12},
  {14.7, 14.5, 11.8},
  {14.4, 14.4, 11.4},
  {14.1, 13.4, 10.4},
  {13.5, 12.4, 9.7},
  {12.6, 12.6, 9.7},
  {12.2, 12.9, 9.6},
  {11.7, 11.1, 7.9},
  {9.9, 9.8, 6.7},
  {9.9, 11, 6.2},
  {11.9, 13.3, 7},
  {14.5, 15.8, 10.1},
  {15.5, 16.9, 12.6},
  {16.6, 17.9, 16.4},
  {17, 19.2, 16.7},
  {16.8, 19.7, 17.6},
  {16.9, 18.8, 17.2},
  {17, 18.3, 15.2},
  {17.3, 18.2, 16.2},
  {16.3, 17.5, 15.9},
  {14.1, 15.7, 13.5},
  {12.3, 13.3, 12.2},
  {12.5, 12.2, 10.9},
  {11.4, 12.1, 9.6},
  {10, 11.1, 9.2},
  {9.3, 10.3, 8.8},
  {8.8, 9.6, 8.7},
  {8.5, 9.1, 7.8},
  {8, 8.7, 7.1},
  {6.5, 7.8, 6.4},
  {6.1, 7.3, 6.1},
  {5.8, 7.5, 5.9},
  {5.7, 7.3, 5.5},
  {6.1, 8.2, 6.2},
  {8.8, 11.2, 8.2},
  {11.8, 13.7, 12.8},
  {13.1, 15, 14.8},
  {14.4, 16.4, 15.2},
  {16.1, 17.9, 15.3},
  {17.1, 18.8, 15.8},
  {17.7, 20.2, 17.1},
  {17.3, 19.2, 16.1},
  {16.7, 17, 15.4},
  {17.3, 19.1, 15.5},
  {15.7, 14.4, 14.2},
  {12.5, 12.3, 10.7},
  {10.6, 12.5, 9.6},
  {9.1, 10.8, 8.4},
  {10.2, 9.9, 7.2},
  {9.1, 9.4, 5.7},
  {8.7, 9.1, 5.4},
  {8.6, 8.7, 4.9},
  {7.7, 8.8, 4.8},
  {7.6, 8, 4.2},
  {7.1, 7.8, 4},
  {7, 7.5, 3.8},
  {6.8, 6.8, 3.6},
  {7.5, 8.2, 4},
  {10.7, 11.2, 6.3},
  {13.2, 13.9, 11},
  {14.2, 15.4, 15.5},
  {15.1, 17, 17},
  {16.6, 19.1, 18.1},
  {17.8, 19.6, 18.8},
  {18.4, 20.7, 19.9},
  {18.9, 21.3, 20.7},
  {19.2, 22.5, 21},
  {19.1, 19.7, 21},
  {16, 15.3, 16.5},
  {14.5, 12.9, 12.1},
  {11.7, 11.4, 10.4},
  {10.7, 10.6, 9.5},
  {10.2, 10.3, 8.5},
  {10.3, 10, 7.9},
  {10, 9.7, 7.4},
  {9.5, 9.1, 6.9},
  {9.2, 9.1, 6.6},
  {9, 8.6, 6},
  {8.7, 8.1, 6},
  {9.2, 7.6, 5.7},
  {8.5, 7.4, 5.7},
  {9, 8.8, 5.8},
  {11.8, 11.2, 7.6},
  {13.9, 13.5, 11.4},
  {14.8, 14.8, 15.9},
  {16.9, 16.4, 18.8},
  {17.8, 18.3, 19.4},
  {18.6, 19.6, 20.1},
  {19, 21.4, 21.1},
  {19.7, 21.7, 21.9},
  {19.3, 22.4, 21.5},
  {19.1, 21.6, 20.8},
  {16.5, 17.7, 19},
  {15.3, 14.8, 16},
  {13, 13.3, 14.1},
  {12.3, 12.7, 12},
  {11.9, 12.2, 11},
  {11.1, 11.6, 10.3},
  {11.1, 11.3, 10},
  {10.9, 10.9, 9.5},
  {10.7, 10.6, 9.1},
  {10.2, 10.4, 8.9},
  {10, 10.1, 8.6},
  {10, 9.8, 8.3},
  {9.7, 9.7, 8.1},
  {10.4, 10.6, 8},
  {13.3, 13.3, 9.5},
  {16.3, 15.5, 14},
  {16.6, 17, 17.5},
  {17.9, 18.8, 19.7},
  {19.1, 20.4, 21.5},
  {20, 21.2, 22.4},
  {21.1, 23, 23.4},
  {21.3, 24.3, 23.7},
  {21, 23.8, 23.3},
  {19.6, 23.3, 23.2},
  {17.8, 19.4, 20.8},
  {16.3, 16.3, 17.8},
  {14.4, 14.7, 16.1},
  {14, 14.9, 14.8},
  {13.6, 14.6, 13.7},
  {13, 14, 13.2},
  {12.9, 13.3, 12.4},
  {12.7, 13.4, 12.4},
  {12.7, 13.2, 12.4},
  {12.9, 12.9, 12.6},
  {12.7, 12.5, 12},
  {12.8, 12.3, 11.4},
  {13.1, 12.4, 11.2},
  {13.8, 13.4, 12.7},
  {16, 16, 14.9},
  {17.4, 16.5, 15.8},
  {19, 18.7, 18},
  {19.3, 19.7, 19.6},
  {20.4, 21.3, 21.8},
  {21.2, 22.4, 23.1},
  {22.1, 23.4, 24.6},
  {22, 24.3, 24},
  {21.9, 24.9, 24.3},
  {20.4, 24.4, 24},
  {19.2, 20.7, 22.2},
  {17.9, 18.2, 19.1},
  {16, 16.5, 17},
  {15.3, 16.1, 16.4},
  {14.9, 15.6, 14.8},
  {14.9, 15.2, 14.4},
  {16, 14.8, 13.8},
  {14.9, 14.5, 13.2},
  {14.5, 14.4, 13},
  {14.1, 14.1, 12.4},
  {13.9, 13.9, 12.4},
  {13.7, 13.7, 11.7},
  {13.6, 13.5, 11.7},
  {14.3, 14.4, 11.9},
  {16.9, 16.6, 13.5},
  {19.2, 19, 18},
  {20, 20.7, 21.1},
  {21.9, 22.1, 24.1},
  {22.2, 23.4, 27},
  {23.2, 24.8, 28.8},
  {24, 26.1, 29.7},
  {25, 27.1, 30.2},
  {24.1, 28, 28.7},
  {23.5, 25.6, 27.6},
  {21.4, 21.9, 25.2},
  {20, 19.7, 21.4},
  {19.7, 18.7, 19.5},
  {18.5, 18.1, 18.2},
  {17.1, 17.5, 16.8},
  {16.3, 17, 15.9},
  {16.1, 16.8, 15.5},
  {15.9, 16.3, 15.4},
  {15.6, 15.8, 14.7},
  {15.3, 15.4, 14.4},
  {15.1, 15.2, 14.2},
  {15.2, 15, 13.8},
  {15.3, 14.7, 13.7},
  {15.7, 15.4, 14.1},
  {18.1, 17.7, 15.1},
  {21.5, 20.4, 18.9},
  {22.7, 22.3, 22.4},
  {23.5, 23.8, 25.1},
  {24.2, 24.9, 27.7},
  {25.2, 26.4, 29.7},
  {26, 27.7, 30.4},
  {26.2, 28.2, 30.5},
  {26.5, 28, 30.3},
  {27.3, 24.9, 29.3},
  {22.4, 21.3, 24.5},
  {19.5, 19.3, 20.3},
  {18.8, 18.5, 18.1},
  {17.8, 18.2, 16.9},
  {17.6, 17.7, 16.2},
  {17.3, 17.3, 15.2},
  {16.6, 16.9, 15},
  {16.6, 16.3, 14.4},
  {17.6, 16.1, 14.3},
  {17.4, 15.6, 13.6},
  {15.7, 15.2, 13},
  {15.1, 14.5, 13.1},
  {15, 14.1, 12.4},
  {15.7, 15, 12.1},
  {18, 17.9, 13.6},
  {21.7, 20.3, 16.5},
  {22.7, 21.6, 21.2},
  {23.5, 23, 24.3},
  {24.4, 24.4, 26.3},
  {24.5, 25.7, 26.5},
  {25.4, 26.8, 27.2},
  {25.6, 27.9, 27.4},
  {25, 27.3, 26.9},
  {24.8, 26, 26.2},
  {22.3, 24.7, 24.4},
  {21.2, 21.8, 21.3},
  {20.8, 19.5, 20},
  {20.9, 19.3, 18.6},
  {20.5, 18.8, 17.5},
  {19.2, 18.3, 16.8},
  {18.8, 18, 16.7},
  {17.5, 18, 16.5},
  {17.2, 17.3, 16.8},
  {17, 17.2, 16.7},
  {17.1, 17.5, 16.3},
  {16.5, 16.8, 16.3},
  {16.8, 16.1, 16},
  {16.9, 16.7, 16.5},
  {18.6, 19.1, 18.1},
  {21, 21.5, 21.3},
  {22.3, 22.8, 22.8},
  {22.9, 23.7, 23.9},
  {23.9, 25.3, 25.1},
  {24.7, 26, 25.9},
  {24.9, 27, 26.8},
  {25, 27.2, 26.8},
  {23.8, 26.6, 25.5},
  {22.1, 25.9, 25.3},
  {21.7, 24, 23.7},
  {20.9, 21.1, 21.6},
  {20.2, 18.8, 19.8},
  {18.6, 18, 18.7},
  {19.5, 17.6, 18.5},
  {19.3, 17.4, 17.8},
  {19, 17, 17.4},
  {17, 16.7, 17.5},
  {17.2, 16.5, 17.4},
  {17.5, 16.6, 16.4},
  {16.7, 16.4, 15.5},
  {16.6, 16.9, 15},
  {16.3, 17.1, 15},
  {16.4, 17.3, 15.1},
  {17.5, 18.6, 16.2},
  {18, 18.9, 16.9},
  {19, 20.6, 18},
  {19.1, 21.2, 20.3},
  {21, 23.4, 23.3},
  {22.2, 24.1, 23.9},
  {22, 23.6, 23.9},
  {22.8, 24.5, 25},
  {23.7, 25.7, 26},
  {23.6, 23.2, 25.2},
  {21.1, 20.9, 20.5},
  {19.4, 21.9, 17.1},
  {19, 20.9, 15.4},
  {18.8, 20.3, 14.3},
  {18.7, 20.4, 13.5},
  {16.8, 18.5, 13},
  {16.5, 16.4, 12.2},
  {15.7, 15.2, 11.4},
  {15.6, 14.5, 10.9},
  {16.1, 14.7, 10.3},
  {15.2, 14.5, 10.2},
  {14.4, 13.1, 10},
  {14.5, 13.4, 9.6},
  {14.2, 13.5, 10},
  {13.6, 15, 10.8},
  {14.2, 17, 15},
  {15.4, 18, 18.7},
  {17, 19.3, 20.4},
  {18.4, 20.4, 21.7},
  {19.2, 21.5, 22.5},
  {19.2, 22.2, 22.8},
  {19.4, 22.8, 23},
  {19.1, 22.9, 22.8},
  {18.6, 22.7, 22.2},
  {16.4, 18.2, 20},
  {13.5, 15.1, 17.9},
  {11.7, 13.6, 15.9},
  {11.5, 12.8, 14.4},
  {11.3, 11.9, 13},
  {11.2, 11.4, 12.4},
  {10.9, 10.8, 11.8},
  {10.5, 10.4, 11.3},
  {10.4, 9.9, 10.7},
  {10.1, 9.4, 10.6},
  {9.9, 9.5, 10.1},
  {9.9, 9.5, 9.8},
  {9.6, 9.6, 9.7},
  {10.1, 10.6, 9.9},
  {12.1, 13.4, 11},
  {16.1, 16.4, 15.6},
  {16.6, 17.4, 18.2},
  {17.4, 18.7, 20.2},
  {18.3, 20.4, 21.9},
  {19.2, 21.5, 22.8},
  {20.2, 22.6, 23.7},
  {20.7, 23.8, 24},
  {20.2, 24.4, 23.9},
  {19.5, 22.5, 23.1},
  {16.7, 18.4, 20.7},
  {14.5, 15.7, 17.6},
  {12.9, 14.8, 16.2},
  {12.7, 13.8, 14.8},
  {12.6, 13, 13.3},
  {12.3, 12.4, 12.7},
  {11.7, 11.9, 11.9},
  {11.5, 11.3, 11.7},
  {11.4, 10.9, 11.2},
  {11.4, 10.9, 10.9},
  {10.9, 10.8, 10.6},
  {10.4, 11, 10.3},
  {10.4, 11, 10.1},
  {10.6, 11.4, 10.1},
  {12.4, 13.6, 11.6},
  {16.6, 16.5, 15.9},
  {17.8, 18, 18.8},
  {18.1, 19.3, 21.2},
  {19.1, 21.1, 23},
  {20.1, 22.4, 23.4},
  {20.8, 23.8, 24.2},
  {21.2, 24.6, 23.4},
  {20, 24.9, 23.8},
  {19.9, 22.3, 21.9},
  {17, 19.4, 19.7},
  {14.6, 17.7, 17.2},
  {13.7, 14.2, 15.8},
  {13.4, 13.2, 13.9},
  {12, 12.1, 12.2},
  {12.5, 11.6, 11.2},
  {13.3, 10.8, 10.1},
  {11.9, 10.7, 9.5},
  {11.3, 9.6, 9.1},
  {10.3, 9.4, 8.2},
  {10.3, 9.2, 8.1},
  {9.8, 8.6, 7.9},
  {9.1, 8.3, 7.4},
  {9.9, 9.2, 7.4},
  {11.9, 12.6, 8.8},
  {15.4, 15.6, 13.1},
  {16.9, 17.3, 17.3},
  {17.8, 18.4, 19.7},
  {18.8, 20.3, 21.3},
  {19.7, 21.6, 22.8},
  {20.7, 22.5, 23.1},
  {20.9, 23.1, 23.1},
  {20.4, 21.9, 23},
  {19, 21.3, 22.4},
  {17, 18.2, 19.7},
  {15.6, 16.9, 16.3},
  {13.3, 17.1, 14.4},
  {12.1, 14.6, 12.5},
  {11.6, 12.7, 11.2},
  {11.7, 12, 10.7},
  {11.8, 11, 10},
  {11.4, 10.4, 9.2},
  {10.8, 9.5, 8.5},
  {9.9, 9.1, 8.1},
  {9.6, 8.6, 7.7},
  {9.3, 8.5, 7.8},
  {9.2, 8.7, 7.3},
  {9.8, 9.1, 7.3},
  {12.4, 12.3, 8.7},
  {15.6, 15.7, 13.4},
  {16.4, 16.8, 16.4},
  {17.7, 18.2, 19.1},
  {18.8, 19.3, 20.1},
  {19.9, 20.8, 21},
  {20, 22.3, 22},
  {20, 22.8, 22},
  {19.3, 22.3, 22},
  {18.9, 21, 21.1},
  {17.1, 18.9, 18.8},
  {16.2, 16.4, 16.3},
  {15.6, 14.9, 14.7},
  {13.2, 13.9, 13.1},
  {12, 13.9, 11.9},
  {12.1, 13.4, 11},
  {13.2, 13, 10.3},
  {12.7, 14, 10.2},
  {13.5, 13.5, 10.6},
  {13.4, 13.6, 10.1},
  {12.8, 12.7, 10},
  {12.8, 12.1, 10},
  {12.9, 12.4, 8.9},
  {13.9, 12.9, 9.6},
  {14.5, 13.3, 12},
  {15.2, 13.6, 12.5},
  {16.3, 14.8, 13.2},
  {16.9, 16.2, 14.6},
  {17.9, 18.4, 16},
  {18.6, 19.5, 17.4},
  {17.5, 19.7, 17.8},
  {17.6, 19.9, 18.3},
  {17.3, 18.2, 18.1},
  {15.7, 17.5, 16.8},
  {14.6, 16.8, 14.6},
  {13.5, 15, 13.3},
  {13.2, 15.4, 12.8},
  {13.5, 14.7, 12.6},
  {13.5, 14.6, 12.8},
  {13, 14.8, 12.7},
  {12.9, 14.1, 12.8},
  {13, 13.6, 12.4},
  {12.5, 13.5, 12.5},
  {12.3, 13.1, 12.3},
  {11.9, 12.9, 11.9},
  {11.8, 12.6, 11.6},
  {11.8, 12.4, 11.4},
  {11.7, 12.4, 11.4},
  {11.9, 12.5, 11.2},
  {12.2, 12.5, 11.9},
  {12.1, 12.8, 12.2},
  {12.5, 13, 12.2},
  {13.7, 13.2, 12.6},
  {14.1, 13.7, 12.5},
  {14, 14.1, 12.9},
  {14.4, 14.6, 13.3},
  {15.6, 14.6, 13.4},
  {16.1, 15.2, 14.1},
  {15.9, 15.3, 14.2},
  {15.5, 14.8, 13.5},
  {15.3, 14.7, 13.2},
  {15.3, 14.9, 13.5},
  {15.8, 15, 13.5},
  {15.3, 15.1, 13.3},
  {13.3, 14.1, 12.8},
  {13.3, 13.7, 11.8},
  {13.2, 14.2, 12},
  {12.4, 13.9, 12},
  {12.3, 12.7, 12.3},
  {12, 11.9, 11},
  {12, 11.4, 10.5},
  {12, 11.6, 10.9},
  {12.6, 13.1, 11.6},
  {13.7, 14.1, 12.7},
  {14.7, 15.2, 14.8},
  {16.1, 15.9, 16},
  {17.9, 18.6, 17.5},
  {18, 19.3, 19},
  {17.7, 19.3, 19},
  {17.6, 20.1, 20.5},
  {17.7, 20.2, 18.8},
  {16.7, 18.6, 16.3},
  {15.2, 15.9, 15},
  {13.9, 15, 14.3},
  {13.6, 14.7, 13.6},
  {13.8, 14.9, 13.3},
  {13.7, 14.3, 13.1},
  {13.5, 14.1, 12.9},
  {13.1, 14.1, 12.5},
  {13.3, 14, 12.2},
  {13.2, 13.8, 12},
  {13, 13.5, 11.6},
  {12.5, 13.5, 11.5},
  {12.3, 13.2, 11.2},
  {12, 13.3, 11.1},
  {12.1, 13.5, 11.1},
  {12.6, 13.1, 11.8},
  {12.3, 12.8, 12.4},
  {12.5, 13.3, 13},
  {13.1, 14.2, 14.5},
  {14.9, 14.9, 16.3},
  {15.9, 16, 16.8},
  {16.1, 15.8, 16.9},
  {15.5, 16, 16.4},
  {15.1, 14.9, 16.4},
  {14.3, 14.8, 15.5},
  {13.8, 14.4, 14.5},
  {12.5, 13.6, 13.3},
  {12.4, 13.1, 12.6},
  {12.1, 12.8, 12.2},
  {11.8, 12.4, 11.9},
  {11.1, 12.2, 11.9},
  {11.1, 11.7, 11.8},
  {11.1, 11.5, 11.4},
  {10.2, 11.8, 10.9},
  {9.7, 12.1, 10.2},
  {9.6, 12.4, 10.2},
  {9.6, 12.3, 10.2},
  {9.7, 12.2, 9.8},
  {10, 12.2, 9.4},
  {10.9, 13.2, 9.9},
  {14.6, 15, 11.8},
  {16.2, 17, 15.8},
  {16.4, 18, 17.6},
  {17.5, 19.5, 18.8},
  {18.3, 19.8, 19},
  {19.3, 20.3, 19.1},
  {19.8, 20.2, 16.3},
  {19, 20.6, 14.9},
  {17, 19.4, 15},
  {15.9, 17.7, 14.3},
  {14.5, 16.2, 13.8},
  {14.2, 14.9, 13.2},
  {14, 14, 13},
  {13.4, 13.8, 12.5},
  {12.5, 13.1, 11.7},
  {11.9, 12.2, 11.4},
  {11.9, 11.7, 10.7},
  {11.5, 11.4, 10.3},
  {11.5, 11.5, 9.6},
  {11.5, 11.8, 9.3},
  {11.2, 11.7, 9.4},
  {11.1, 11.7, 9.5},
  {11.6, 12.4, 10},
  {13.6, 12.9, 10.9},
  {15.9, 14.4, 13},
  {16.2, 16.4, 14.8},
  {17, 17.8, 18.8},
  {18.6, 20.2, 19.6},
  {19.5, 20.1, 19.4},
  {19.9, 21.7, 20.7},
  {19.7, 19.5, 22},
  {19.6, 21.2, 19.7},
  {19.1, 17, 19.9},
  {16.6, 15.9, 16.6},
  {14.6, 14.5, 15.1},
  {13.3, 14.1, 14.4},
  {14, 12.9, 12.8},
  {14, 12.2, 11},
  {13.4, 12.2, 10.4},
  {13.1, 12.5, 9.8},
  {12.5, 12.1, 9.9},
  {12, 11.7, 9.9},
  {11.4, 11.2, 8.9},
  {10.8, 10.3, 8.6},
  {10.4, 9.7, 7.9},
  {10.3, 9.4, 7.5},
  {10.1, 9.6, 7.5},
  {11.1, 12.4, 8.7},
  {15.3, 15.5, 12.4},
  {16.3, 16.9, 15.3},
  {17.1, 18.2, 18.6},
  {18.3, 18.9, 20.1},
  {19.2, 20, 20.7},
  {19.9, 21, 21.2},
  {20, 20.1, 21.4},
  {18.6, 20, 21.1},
  {17.7, 18.1, 20.3},
  {16.5, 15.7, 17.4},
  {15.2, 14.3, 14.3},
  {13.7, 13.5, 12.9},
  {13.2, 13.4, 11.8},
  {12.8, 12.9, 11.3},
  {13.4, 12.5, 11},
  {14.2, 12.4, 10.5},
  {14.4, 12.8, 9.9},
  {14.2, 13.2, 9.9},
  {13.9, 13.3, 10.4},
  {14, 12.5, 10.8},
  {13.6, 12.8, 10.9},
  {13.4, 12.6, 11.3},
  {13.5, 12.8, 10.8},
  {14.2, 13.6, 11},
  {15.2, 15.3, 13.4},
  {16.1, 17.7, 17.2},
  {17.3, 18.4, 19.5},
  {18.2, 20, 19.9},
  {19.2, 20.9, 20.6},
  {19.8, 21.8, 20.9},
  {19.6, 22.6, 20.9},
  {19.5, 21.5, 21},
  {18.3, 17.8, 20.5},
  {16.5, 16.1, 18.3},
  {15.9, 14.8, 15.4},
  {15.5, 13.8, 14.8},
  {15.1, 13.5, 14.7},
  {15.2, 13.4, 14.6},
  {14.6, 13.4, 14.2},
  {14.5, 13.2, 14},
  {14.9, 13.4, 13.8},
  {14.8, 13.7, 13.3},
  {14.6, 14, 12.8},
  {14.4, 13.9, 12.7},
  {13.5, 13.7, 12.6},
  {12.9, 12.9, 12},
  {12.4, 12.5, 11.7},
  {14, 13.8, 11.6},
  {16, 16.4, 14.5},
  {17.5, 17.7, 17.5},
  {18.6, 19.3, 19.5},
  {19.1, 20.6, 20.6},
  {19.7, 21.8, 21.3},
  {20.1, 22.4, 22.2},
  {20, 23.2, 22.2},
  {18.6, 22.8, 21.7},
  {17.7, 18.8, 20.7},
  {17.1, 16.5, 18.6},
  {16.8, 15, 16.3},
  {16.9, 14.4, 14.9},
  {16.1, 14.3, 14},
  {15.9, 14, 14.7},
  {16.1, 15.1, 14.3},
  {16.2, 15.7, 14.2},
  {16, 15.8, 14.3},
  {15.9, 15.7, 14.4},
  {15.7, 15.6, 14.4},
  {15.7, 15.6, 14.2},
  {15.6, 15.5, 14.1},
  {15.5, 15.5, 14},
  {15.2, 15.6, 14},
  {15.1, 15.8, 14.6},
  {14.9, 16.4, 15.2},
  {15, 17.4, 15.9},
  {15.9, 18.2, 16.9},
  {16.1, 18.7, 18.2},
  {16.6, 19.3, 19.2},
  {17.4, 19.9, 20.3},
  {16.7, 20, 19.7},
  {16.4, 19.6, 19.2},
  {16.2, 18.8, 18.3},
  {15.3, 17.5, 16.9},
  {14.5, 15.1, 16.1},
  {13.8, 14.9, 15.6},
  {12.3, 14.4, 15},
  {11.7, 13.8, 14.6},
  {11.7, 13.1, 14.3},
  {11.9, 13.4, 14.1},
  {11.7, 13.1, 12.7},
  {10.9, 11, 12.9},
  {11.3, 11.7, 12.9},
  {9.7, 11.7, 12},
  {9.4, 10, 11.4},
  {9.8, 9.7, 11.7},
  {11.6, 9.8, 11.9},
  {11.6, 12.9, 13.3},
  {14.2, 14.8, 15.3},
  {15.4, 16.2, 16.4},
  {16.2, 17.5, 17.6},
  {17, 18.7, 18.5},
  {17.5, 19.8, 17.6},
  {17.7, 19.8, 18.1},
  {17.1, 18.9, 18.3},
  {15.6, 19, 17.9},
  {14.5, 17.5, 16.6},
  {14.2, 15.3, 15.9},
  {13.6, 13.8, 15.3},
  {13, 12.9, 13.8},
  {12.1, 12.4, 12.8},
  {11.6, 12.2, 11.7},
  {12, 11.8, 11},
  {12.3, 12.2, 10.9},
  {11.8, 12.3, 10.6},
  {11.5, 12, 10.1},
  {12, 11.6, 10.1},
  {11.9, 12, 9.8},
  {12.5, 11.6, 8.9},
  {12.4, 11.2, 8.3},
  {12.6, 11.8, 8.7},
  {13, 12.3, 10.4},
  {13.3, 13.6, 13.1},
  {13.5, 14.4, 13.9},
  {13.4, 15.4, 14.7},
  {13.2, 15.8, 15.9},
  {13.1, 16.2, 15.9},
  {13.8, 16.2, 15.9},
  {13.9, 15.6, 15.2},
  {13.7, 15.5, 14.9},
  {13.1, 15.2, 14.4},
  {12.9, 14.3, 13.4},
  {12.9, 14.2, 12.4},
  {12.7, 14.1, 11.9},
  {12.1, 13.4, 11.6},
  {11.7, 13.5, 11.2},
  {12.1, 13.8, 11},
  {12.4, 13.5, 10.9},
  {12.4, 12.9, 10.5},
  {12.6, 12.5, 10.3},
  {12.7, 11.9, 10.3},
  {12.5, 11.6, 10.2},
  {12.5, 11.5, 10},
  {12.7, 11.6, 9.8},
  {12.3, 10.9, 9.4},
  {12.9, 12, 10.5},
  {14.5, 14.2, 12},
  {14, 16, 13.8},
  {14.8, 16.8, 15.6},
  {16.4, 17.5, 16.8},
  {17.2, 17.9, 18.8},
  {18, 19.6, 20},
  {18.1, 21.1, 19.9},
  {18.2, 20.8, 19.8},
  {17.5, 20.1, 18.8},
  {15.3, 16.8, 16.1},
  {14.1, 14.7, 14.2},
  {13.5, 13.4, 12.6},
  {12.8, 12.3, 11.5},
  {13.4, 11.6, 11.1},
  {14.4, 11.6, 11.5},
  {13.7, 11.8, 11.6},
  {13, 12.2, 11.5},
  {13.5, 12.3, 10.8},
  {13.8, 11.6, 9.9},
  {13.4, 10.5, 9.1},
  {12.6, 10.8, 8.4},
  {10.7, 10.6, 8},
  {10.8, 10.3, 8.2},
  {11.5, 13, 9},
  {15.6, 16.2, 11.4},
  {16.1, 17.3, 14.9},
  {17.1, 18.5, 18.2},
  {18, 19.9, 19.6},
  {19.1, 21, 18.3},
  {19.6, 21.2, 21.6},
  {19.5, 18.2, 20},
  {18.9, 15.8, 19.9},
  {17.6, 16.1, 16.6},
  {15.9, 13.9, 15.2},
  {13.5, 13.4, 14},
  {12.5, 12.4, 12.7},
  {12.1, 12.9, 12.3},
  {12.8, 13.5, 12.1},
  {12.6, 13.6, 12.1},
  {13, 13.3, 11.3},
  {12.9, 12.5, 10.8},
  {12, 12.1, 10.7},
  {13.3, 12.1, 10.9},
  {13.1, 12.1, 10},
  {11.4, 11.8, 9.7},
  {10.9, 10.7, 9.4},
  {11, 11, 9.2},
  {12.2, 13.7, 9.7},
  {15.3, 15.3, 12.5},
  {16.6, 17.1, 15.9},
  {17, 17.6, 18.5},
  {17.8, 19.1, 19.4},
  {18.2, 19.8, 19.4},
  {18.5, 20.7, 20.3},
  {18.5, 21.6, 20.5},
  {18.2, 18.6, 20.7},
  {17, 16.6, 19.4},
  {15.4, 14.6, 16.8},
  {14.3, 13.4, 14.7},
  {12.6, 12.7, 13.3},
  {12.4, 12.4, 12.4},
  {12.1, 11.9, 11.5},
  {11.8, 11.7, 11.3},
  {11.7, 11.5, 11},
  {11.2, 11.4, 10.4},
  {11.3, 11.6, 10},
  {11.3, 11, 10.1},
  {11.2, 10.5, 9.5},
  {11.2, 10.5, 8.8},
  {11.3, 10.7, 8.8},
  {11.3, 10.6, 9.6},
  {12.5, 11.6, 10.7},
  {14.9, 15, 12.7},
  {15.6, 16.6, 16},
  {17, 17.8, 18.3},
  {18, 18.8, 17.9},
  {18.5, 20.1, 18.9},
  {18.6, 20.8, 18.9},
  {17.9, 21, 18.1},
  {17.3, 20.7, 16.7},
  {_, 17.6, 16.5},
  {16.7, 15.9, 15.4},
  {14.6, 13.7, 14},
  {14.5, 12.9, 13.2},
  {12.8, 12.6, 12.6},
  {12.4, 12.1, 12.1},
  {12, 11.9, 12.2},
  {11.5, 11.8, 11.9},
  {11.6, 11.5, 11.1},
  {11.6, 11.7, 11.1},
  {11.7, 11.4, 11},
  {11.4, 11.5, 10.9},
  {10.8, 11.1, 9.5},
  {11, 11, 9},
  {11.5, 11.1, 9},
  {12.6, 11.9, 10.2},
  {14.4, 14.3, 13},
  {16.5, 16.4, 15.1},
  {17.2, 17.5, 17.4},
  {17.8, 19, 16.7},
  {18.1, 19.4, 19.4},
  {18.1, 20, 20.1},
  {18.2, 20, 19.8},
  {16.3, 19.3, 19.3},
  {15.8, 17.9, 17.7},
  {15.4, 15.9, 16.3},
  {14.9, 14.7, 14.6},
  {14.1, 14.8, 13.7},
  {13.3, 14.7, 13.2},
  {13.9, 13.7, 12.9},
  {12.6, 13.4, 13},
  {12.2, 12.6, 12.2},
  {12.5, 12.2, 11.8},
  {12.2, 12.2, 11.8},
  {11.7, 12.1, 11.1},
  {11.8, 11.9, 11.4},
  {12.6, 12.1, 11.4},
  {13, 12, 11},
  {13.1, 12.5, 10.6},
  {13.5, 13.3, 11.4},
  {13.8, 14.3, 15.1},
  {14.3, 14.9, 16.2},
  {15.3, 15.8, 16.6},
  {16, 17.6, 18.7},
  {16.3, 19, 19.9},
  {16.1, 18.8, 19.5},
  {16.1, 18.8, 18.9},
  {15.8, 18.5, 18.3},
  {15.2, 17.7, 17.6},
  {15, 16.7, 15.8},
  {15.2, 16, 14.6},
  {15.3, 15.7, 14.3},
  {15.3, 15.6, 13.9},
  {15.4, 15.7, 13.9},
  {15.5, 15.6, 13.8},
  {15.2, 15.4, 13.8},
  {14.7, 15.2, 13.7},
  {14.5, 15.5, 13.5},
  {14.5, 15.3, 13.5},
  {14.5, 15.3, 13.4},
  {14.5, 15.1, 13.5},
  {14.3, 15.1, 13.3},
  {14.1, 15.2, 13.3},
  {14.4, 15.5, 13.6},
  {14.8, 16.1, 14.5},
  {15.5, 16.3, 15.5},
  {16.5, 16.6, 16.1},
  {17.3, 17.6, 17.8},
  {17.2, 19, 17.6},
  {17.8, 19.9, 18.7},
  {18.8, 20.8, 19.1},
  {18.1, 21, 18.7},
  {17.6, 19.7, 18.3},
  {16.5, 17.8, 16.5},
  {15.9, 15.8, 15.4},
  {15.3, 14.8, 14.6},
  {14.8, 14, 13.7},
  {15.5, 13.9, 12.2},
  {15.3, 13.8, 11.7},
  {15.2, 13.9, 11.8},
  {14.9, 14, 12.1},
  {14.9, 13.7, 12.1},
  {14.9, 13.4, 11.9},
  {14.9, 13.7, 11.1},
  {14.7, 14, 10.1},
  {14.8, 14.2, 9.9},
  {14.8, 14, 10.4},
  {14.9, 14.9, 12.5},
  {14.9, 15, 13.2},
  {15, 15.5, 13.3},
  {15.2, 15.4, 14},
  {15.1, 15.4, 14.3},
  {15, 15.2, 14.3},
  {15.3, 15.3, 14.4},
  {15.7, 15.4, 14.5},
  {16.1, 15.4, 14.9},
  {16.7, 15.3, 14.8},
  {16.9, 16.3, 16.3},
  {17.3, 16.6, 17.2},
  {17.2, 17.8, 17.2},
  {16.8, 16.1, 15.2},
  {17.3, 16.3, 15.8},
  {17.2, 15.8, 17.1},
  {17, 16.1, 17.3},
  {16.8, 16.2, 16.5},
  {16, 15.9, 14.5},
  {15.9, 16, 13.7},
  {14.8, 16, 13},
  {14, 14.2, 12.8},
  {12.9, 13.3, 12.6},
  {13.2, 13.3, 12.2},
  {13.5, 12.5, 12.1},
  {13.4, 13.1, 11.5},
  {13.3, 13.8, 11.9},
  {13.2, 15.2, 13.1},
  {14.1, 15.8, 15.4},
  {15, 15.6, 16.2},
  {15.8, 15.3, 14.8},
  {14.6, 14.1, 13.2},
  {14.1, 13.2, 11.6},
  {11.9, 12, 10.3},
  {9.9, 10.5, 9.4},
  {8, 9, 7.5},
  {7.1, 7.7, 6.5},
  {6.4, 7.3, 6.1},
  {6, 7.3, 5.4},
  {5.6, 7.3, 5.1},
  {5.2, 7, 5.4},
  {4.5, 6.5, 5.5},
  {4.4, 6.5, 5},
  {4.2, 7.3, 4.6},
  {4.2, 6.7, 4.4},
  {4.1, 5.9, 4.1},
  {4.1, 4.9, 4.4},
  {3.9, 4.9, 4.1},
  {5, 5.8, 5.5},
  {8.4, 7.1, 7.8},
  {10.2, 9.3, 10.2},
  {11.1, 12.4, 12.4},
  {12.4, 14.3, 14.2},
  {13.8, 15.5, 15.4},
  {14.7, 17, 16.5},
  {14.9, 17, 16.7},
  {14.4, 14.5, 16.8},
  {13.3, 10.9, 14.2},
  {11.3, 8.9, 10.1},
  {10.8, 8, 8.5},
  {10.6, 7.8, 7.3},
  {8.4, 7.3, 6.1},
  {7.6, 6.9, 5.3},
  {7.4, 6.7, 4.9},
  {7.8, 6.6, 4.5},
  {7.3, 6.3, 4.3},
  {6.7, 6.1, 4},
  {6.5, 5.7, 3.6},
  {6.4, 5.3, 3.5},
  {6.1, 4.9, 3.4},
  {7.1, 4.5, 3.1},
  {6.7, 4.5, 2.9},
  {7.5, 6.7, 4.1},
  {9.1, 8.1, 7.1},
  {10.4, 10.1, 9.5},
  {11.6, 11.6, 12.3},
  {12.2, 13.1, 14.2},
  {13.3, 14, 14.9},
  {14.1, 15.7, 15.7},
  {14.3, 16.5, 16},
  {13.7, 14.5, 15.6},
  {12.2, 10.8, 14.1},
  {10.5, 9.6, 11},
  {8.7, 8.7, 9.2},
  {8.6, 8.2, 7.6},
  {9.1, 7.8, 6.6},
  {8.2, 7.5, 6.4},
  {7.9, 7.3, 5.9},
  {8.6, 7.3, 5.5},
  {8.5, 7.2, 5.1},
  {8.8, 7.1, 5},
  {8.1, 7.1, 4.9},
  {7.7, 6.9, 4.9},
  {7.7, 6.6, 4.9},
  {7.6, 6.9, 5.3},
  {7.2, 7.1, 5.6},
  {8.3, 7.8, 5.7},
  {9.6, 9.7, 8.9},
  {10.1, 11.1, 10.1},
  {10.3, 10.8, 12.3},
  {10.7, 10.1, 11.8},
  {10.4, 10.7, 11.5},
  {11, 11.5, 11.7},
  {11.2, 13.2, 12.9},
  {12, 12.9, 13.5},
  {11.9, 10.9, 12.7},
  {9, 9, 10.4},
  {8, 8.3, 8.5},
  {7.7, 8.1, 7.6},
  {7.8, 7.7, 6.9},
  {8.8, 8.8, 5.9},
  {9.1, 10.7, 5.4},
  {8.3, 10.5, 5.2},
  {8.1, 9.2, 4.7},
  {8.2, 9, 4.3},
  {6.7, 8.6, 4.2},
  {6, 8.5, 3.8},
  {5.8, 6.9, 3.8},
  {5.5, 6.3, 3.6},
  {6, 5.6, 3.2},
  {6.1, 7.5, 3.2},
  {10, 10.7, 6.2},
  {12.5, 12.1, 8.8},
  {13.5, 13.3, 12.1},
  {14.4, 14.7, 14.7},
  {15, 15.6, 15.9},
  {15.6, 17.2, 18.1},
  {15.6, 16.9, 17.5},
  {15.2, 14.5, 17.1},
  {14.2, 10.3, 14.9},
  {10.2, 9.1, 9.9},
  {9.5, 8.6, 8.2},
  {9.5, 8.3, 7.2},
  {8.5, 8.2, 6.5},
  {8, 7.8, 6.2},
  {8.2, 7.5, 6},
  {7.4, 6.9, 5.5},
  {7.5, 6.8, 4.7},
  {8.1, 6.7, 4.2},
  {7.8, 6.3, 3.5},
  {7.1, 5.9, 3.2},
  {6.1, 5.4, 3.4},
  {5.9, 5.2, 2.8},
  {5.9, 5, 2.6},
  {6.5, 6.9, 3.2},
  {9.7, 10.2, 7.1},
  {12.5, 11.6, 9.5},
  {13.7, 12.8, 12.7},
  {14.9, 14.6, 16.3},
  {15.6, 16.1, 17.7},
  {16, 16.9, 19.1},
  {16.5, 18.6, 19.8},
  {16.6, 16.5, 18.8},
  {15.1, 11.6, 15.7},
  {11.4, 10.5, 11.4},
  {10.1, 9.6, 10},
  {9.3, 9.2, 9.4},
  {8.9, 8.7, 8.3},
  {9.1, 8.5, 7.8},
  {9.3, 8.2, 7.6},
  {9.1, 7.9, 7.3},
  {8.9, 7.5, 6.6},
  {8.3, 7.3, 6.9},
  {8, 6.8, 6.5},
  {7.6, 6.9, 6.7},
  {7.8, 6.5, 6},
  {7, 6.4, 5.9},
  {7.4, 6.3, 5.3},
  {7.9, 8.1, 5.4},
  {12.1, 12.1, 9.3},
  {14.3, 13.6, 11.6},
  {15.4, 15.2, 14.3},
  {17.1, 16.6, 17.6},
  {18.1, 17.4, 19.4},
  {18.3, 18.3, 20.4},
  {18.5, 19.6, 20.5},
  {18, 16.1, 20.1},
  {15.7, 11.7, 17.4},
  {12, 10.7, 12.4},
  {10.6, 9.9, 10.8},
  {10.3, 9.7, 9.7},
  {10.6, 9.3, 8.7},
  {10, 9.1, 8},
  {9.8, 8.4, 7.9},
  {9.5, 8.1, 7.3},
  {9, 7.8, 6.7},
  {8.3, 7.4, 7},
  {8.1, 7.2, 6.5},
  {8, 6.7, 5.6},
  {7.7, 6.3, 5.5},
  {7.4, 6.3, 5.3},
  {7.3, 6.1, 5.2},
  {7.8, 7.9, 5.7},
  {12.1, 11.9, 9.1},
  {14.5, 13, 11.8},
  {15.3, 14.3, 14.2},
  {16.8, 15.4, 17.3},
  {16.7, 16.9, 18.6},
  {17.3, 17.8, 19.4},
  {17.5, 18.4, 19.4},
  {15.7, 15.1, 18.8},
  {14.6, 11.3, 16.3},
  {12.3, 10.7, 12.3},
  {9.8, 9.9, 10.4},
  {9, 9.4, 8.6},
  {8.2, 8.4, 8},
  {8.3, 8.1, 7.1},
  {8.2, 7.7, 6.7},
  {8.2, 7.7, 6.3},
  {7.9, 7.3, 6.1},
  {7.5, 6.9, 5.7},
  {7.2, 6.8, 5.5},
  {7.1, 7, 5.2},
  {7, 6.9, 5.1},
  {6.8, 6.6, 5.1},
  {6.8, 6.5, 5},
  {7.4, 7.8, 5.2},
  {10.8, 11, 8.1},
  {13.1, 12.4, 10.7},
  {13.6, 13.9, 14.3},
  {14.8, 15.1, 17},
  {15.4, 15.7, 17.8},
  {15.4, 16.7, 19.4},
  {15.5, 18.1, 18.5},
  {15.1, 16.8, 18.4},
  {14.2, 12.2, 16.3},
  {10.6, 10.6, 12.5},
  {9.7, 10, 11},
  {9.3, 9.6, 9.8},
  {9.3, 9.2, 9},
  {9, 9.1, 8.7},
  {9.3, 8.9, 8.2},
  {9.1, 8.8, 7.7},
  {9, 8.6, 7.4},
  {8.8, 8.8, 7.3},
  {8.8, 8.1, 6.9},
  {8.8, 8, 6.7},
  {9.2, 7.8, 6.4},
  {8.8, 7.6, 6.8},
  {9, 7.9, 7.1},
  {9.4, 8.9, 7.8},
  {12.5, 12.9, 9.6},
  {14.4, 14.1, 12.2},
  {16.1, 14.9, 15.8},
  {17.2, 16.1, 17.8},
  {18.6, 17.8, 19.6},
  {18.4, 18.4, 17.4},
  {18.6, 20.4, 17.9},
  {17.5, 19.7, 15.8},
  {16.3, 16.2, 15.2},
  {13.3, 13.9, 13.1},
  {11.6, 11.8, 12.4},
  {11.3, 10.7, 11.4},
  {10.8, 10.5, 11},
  {10.4, 10.1, 10.3},
  {9.9, 10.7, 9.2},
  {9.6, 10.5, 8.4},
  {9.9, 9.8, 7.9},
  {9.8, 9.7, 7.4},
  {9.2, 9.4, 7},
  {8.5, 9.3, 6.4},
  {8.5, 9.3, 6.8},
  {8.5, 8.3, 6.6},
  {8.8, 9, 6.5},
  {10.4, 9.7, 6.7},
  {11.8, 10.6, 8.2},
  {12.2, 11.7, 10.1},
  {12.4, 12.8, 11.3},
  {12.5, 13, 11.8},
  {12.1, 13.3, 12.5},
  {12, 12.9, 12.4},
  {11.8, 12.7, 11.7},
  {11.6, 12.4, 11.3},
  {11.5, 12.4, 11},
  {10.6, 11.8, 10.7},
  {10, 11.4, 10.2},
  {9.8, 11.1, 9.6},
  {10.5, 11.6, 9.3},
  {10.7, 12.4, 9.1},
  {10.4, 12.4, 9},
  {10.2, 12.2, 9},
  {10, 12.1, 9},
  {9.7, 11.7, 8.8},
  {9.4, 11.6, 8.3},
  {9.2, 10.5, 7.9},
  {8.2, 8.1, 7.4},
  {7.2, 8, 6.8},
  {6.9, 6.7, 6.1},
  {7.8, 7.5, 5.7},
  {10.3, 11.4, 6},
  {12.4, 12.8, 8.5},
  {12.2, 13.7, 11.3},
  {13.4, 14.5, 12.8},
  {14.2, 15.5, 13.8},
  {14.8, 16.1, 15},
  {15.3, 16.5, 15.2},
  {14.7, 12.5, 15.1},
  {13.2, 9.4, 12.8},
  {9.8, 8.6, 8.9},
  {8.2, 8.3, 7.6},
  {7.3, 8, 6.8},
  {7.1, 7.5, 6.2},
  {7.5, 7.3, 5.6},
  {7.3, 7, 5.1},
  {6.9, 6.6, 4.8},
  {6.2, 6.7, 4.5},
  {6.2, 6.1, 4.3},
  {5.9, 5.8, 3.8},
  {5.9, 5.1, 3.8},
  {5.8, 5, 3.6},
  {5.7, 4.7, 3.3},
  {5.2, 4.6, 3.2},
  {5.7, 5.7, 3.4},
  {9.7, 9.5, 5.9},
  {12, 10.9, 8.8},
  {13.4, 12.1, 11.2},
  {14.5, 13.4, 14.1},
  {14.4, 15, 16.4},
  {14.7, 15.7, 17},
  {15.2, 15.9, 17},
  {12.9, 13.9, 16.2},
  {11.5, 12.2, 14.1},
  {9.8, 11.7, 10.3},
  {8.2, 11.2, 8.7},
  {9.1, 10.6, 6.6},
  {9.4, 8.1, 5.9},
  {9.3, 8.4, 6.8},
  {9.2, 10.4, 7.2},
  {9.1, 9.6, 7.4},
  {8.8, 8.8, 7.6},
  {8.4, 8.1, 7.4},
  {8.1, 6.8, 7.3},
  {7.9, 6.4, 7.2},
  {7.4, 6, 7.1},
  {7, 5.5, 7},
  {5.2, 5.5, 6.9},
  {5.7, 5.8, 7.4},
  {8, 8, 8.2},
  {8.4, 9.4, 9.4},
  {9.3, 10.8, 10.6},
  {11, 12.8, 13.1},
  {12, 13.5, 13.8},
  {12.4, 13.6, 13.7},
  {12.5, 12.9, 13.5},
  {11.5, 10.1, 12.8},
  {10.3, 8.6, 11.6},
  {6.9, 7.6, 8.8},
  {5.8, 6.5, 7.1},
  {5.3, 6.1, 6.8},
  {4.9, 5.9, 7.8},
  {4.8, 5.3, 7.7},
  {4.6, 5.2, 7.7},
  {4.5, 5, 7.9},
  {4.3, 4.7, 7.7},
  {4.2, 4.8, 7.8},
  {4, 5.7, 7.7},
  {3.9, 7.5, 6.6},
  {4, 7.5, 6.4},
  {4, 7, 6.3},
  {4.2, 6.9, 5.8},
  {6.1, 7.2, 5.5},
  {8.6, 7.9, 5.6},
  {9.7, 9, 8.2},
  {10.5, 9.8, 10.1},
  {11.3, 11.2, 10.8},
  {11.5, 12.8, 12.4},
  {11.8, 13.2, 13.7},
  {12.4, 13.7, 13.3},
  {10.6, 13.6, 12.5},
  {9.2, 11.5, 11.4},
  {7.7, 9.9, 9},
  {6.6, 8.7, 7.6},
  {6.7, 9.2, 6.1},
  {6.5, 9.8, 5.6},
  {6.2, 9.3, 4.9},
  {6, 9.3, 4.9},
  {6.1, 8.5, 4.4},
  {5.7, 7.8, 4.5},
  {6.4, 7.9, 4.4},
  {7, 8, 4.9},
  {7.1, 8.1, 4.5},
  {6.9, 8.1, 3.7},
  {5.8, 8.1, 3.5},
  {5.6, 8.1, 4},
  {7, 8.6, 4.3},
  {7.7, 8.8, 6.1},
  {8.1, 9.1, 8},
  {8.5, 9.5, 9.6},
  {9.4, 9.9, 11.4},
  {10, 10.6, 12.4},
  {10.9, 11.1, 13},
  {10.4, 11.7, 12.9},
  {10.1, 11.8, 11.9},
  {9.4, 11.3, 10.6},
  {9, 10.5, 9.6},
  {9.1, 10, 8.9},
  {9.3, 10, 8.6},
  {9.3, 10.1, 8.4},
  {9, 10.5, 8.1},
  {8.7, 10.5, 7.7},
  {8.6, 10, 7.6},
  {7.9, 9.1, 7.8},
  {7.4, 8.7, 7.1},
  {7, 8.5, 6.9},
  {6.9, 8.4, 6.7},
  {6.8, 8.1, 6.6},
  {6.8, 7.8, 6.5},
  {6.9, 7.7, 6.6},
  {7, 8.2, 6.8},
  {7.3, 8.5, 7.2},
  {7.4, 8.8, 7.9},
  {7.7, 9, 9},
  {8.6, 9.6, 9.7},
  {9.6, 10.3, 10.7},
  {10.6, 10.8, 12.6},
  {10.7, 12, 12.3},
  {10.5, 12.1, 11.4},
  {10.1, 11.3, 10.9},
  {8.5, 10.6, 10.3},
  {7.5, 10.1, 9.9},
  {8.3, 9.9, 9.6},
  {8.4, 9.5, 9.3},
  {8.8, 9.3, 9},
  {9.1, 9.7, 8.8},
  {8.8, 9.9, 8.6},
  {8.6, 9.7, 8.7},
  {8.6, 9.5, 8.5},
  {8.5, 9, 8.4},
  {8.6, 8.9, 7.7},
  {8.6, 9.2, 7.3},
  {8.6, 9.5, 6.6},
  {8.7, 9.9, 7},
  {8.8, 9.8, 7.7},
  {8.9, 9.8, 8.5},
  {9.2, 10.2, 9},
  {9.5, 10.6, 9.7},
  {10.2, 10.9, 10.9},
  {10.1, 11.3, 11.1},
  {9.9, 11.9, 11.3},
  {10.4, 12.4, 11.7},
  {10.5, 12.3, 11.9},
  {10.2, 12.1, 11.4},
  {8.6, 10.5, 10.7},
  {8.3, 10, 10.2},
  {7.8, 9.9, 9.8},
  {7.4, 9.6, 9.8},
  {8.3, 9.1, 9.8},
  {8.3, 9.7, 9.6},
  {7.6, 8.9, 9.7},
  {7.5, 9.5, 9.4},
  {7.4, 9.8, 8.9},
  {7.2, 9.3, 8.6},
  {7.1, 9.3, 8.6},
  {7, 8.9, 7.8},
  {7.2, 9.5, 7.1},
  {8.3, 9.5, 6.5},
  {9.1, 9.9, 6.8},
  {10.1, 10.3, 8.9},
  {10.5, 11.1, 11.4},
  {11.3, 11.6, 13},
  {11.9, 12.9, 14.6},
  {13.5, 14.3, 14.9},
  {13.1, 15.2, 16.1},
  {13.7, 15.3, 16.2},
  {13.2, 14.7, 15.3},
  {12, 13.8, 13.1},
  {9.9, 13, 11.1},
  {9.1, 12.2, 9.6},
  {10.3, 12.2, 8.4},
  {10.6, 11.9, 8.9},
  {10.5, 12.3, 8.6},
  {10.5, 12.5, 7.9},
  {9.6, 11.8, 7.9},
  {9.4, 11.8, 7.9},
  {10.1, 11.5, 8},
  {10.2, 11.5, 8},
  {10.3, 11.4, 7.5},
  {10.2, 11.1, 7.6},
  {10, 10.9, 7.3},
  {10, 10.9, 7.4},
  {10.3, 11, 7.6},
  {10.8, 11.2, 9.1},
  {11, 11.6, 10.3},
  {11.1, 11.7, 11.3},
  {11.1, 11.5, 12.4},
  {11.2, 11.3, 11.8},
  {11.5, 11.5, 11.7},
  {11.6, 11.6, 11.4},
  {11.5, 11.6, 11.3},
  {11.5, 11.5, 11},
  {11.7, 11.5, 10.5},
  {11.9, 11.8, 10.5},
  {11.9, 12, 10.3},
  {12, 12.3, 10.3},
  {12.2, 12.5, 10.2},
  {12.2, 12.8, 10.4},
  {12.9, 12.9, 10.5},
  {13.8, 12.7, 10.5},
  {14, 13, 11.3},
  {13.8, 13.3, 11.5},
  {13.6, 13.6, 11.7},
  {13.4, 14, 11.8},
  {13.3, 13.9, 11.8},
  {13.5, 14, 11.8},
  {13.7, 14.1, 11.7},
  {14.3, 14.6, 11.8},
  {14.7, 15, 12.5},
  {15.2, 15.7, 13.2},
  {15.9, 16.8, 13.5},
  {16.4, 15.6, 13.7},
  {16.4, 17, 14.9},
  {17, 18.2, 15.6},
  {16.6, 17.8, 16.3},
  {15.8, 16.7, 14.1},
  {14.5, 14.3, 11.1},
  {14, 14, 10.1},
  {14, 13.7, 9.4},
  {13.3, 13.1, 8.8},
  {12.5, 12.1, 8.7},
  {11.1, 11.6, 8.2},
  {9.5, 11.4, 8},
  {9.4, 11.5, 7.7},
  {9, 11, 7.2},
  {9.6, 10.4, 6.5},
  {8.9, 9.6, 6},
  {9.2, 9.6, _},
  {8.6, 9.9, 5.6},
  {8.6, 9.5, 5.1},
  {8.7, 9.2, 5.1},
  {10.7, 9.7, 8.5},
  {13.9, 10.4, 8.9},
  {14.6, 13.2, 9.8},
  {15.6, 14.8, 12.6},
  {16.1, 16.1, 15.4},
  {16.3, 16.5, 18},
  {16.7, 17.7, 18.9},
  {15.9, 16.4, 18.4},
  {13.6, 15.6, 17.5},
  {12.2, 13.7, 16.3},
  {10.7, 13, 14.3},
  {10.1, 12.1, 12.8},
  {10, 12.5, 11.8},
  {9.6, 12.8, 10.8},
  {9.5, 12.3, 9.9},
  {9.4, 11.8, 9.3},
  {9.4, 11.6, 8.7},
  {9, 11.4, 8.4},
  {8.8, 11.1, 8},
  {8.8, 10.9, 8.2},
  {8.7, 10.9, 8.1},
  {8.6, 10.5, 7.7},
  {8.4, 10.6, 8.2},
  {8.8, 10.6, 8.7},
  {10.6, 11.3, 9.2},
  {13.5, 11.3, 9.3},
  {15.1, 14.9, 9.7},
  {15.7, 16, 12.1},
  {16.5, 17.1, 16},
  {16.8, 18.1, 19.2},
  {16.9, 18.1, 20.3},
  {15.5, 17.9, 18.6},
  {13.7, 16.1, 17.4},
  {11.9, 13.7, 15.3},
  {11, 12.8, 13.2},
  {11.5, 12.7, 12},
  {11.6, 12.4, 11.8},
  {11.6, 12.2, 11.5},
  {11, 12.2, 10.8},
  {10, 11.5, 10.3},
  {10, 11.2, 10},
  {10.4, 11.2, 9.3},
  {10, 11.7, 9},
  {9.4, 11.6, 8.7},
  {9.2, 11.5, 9.2},
  {8.8, 11.2, 9.6},
  {8.4, 10.9, 9.6},
  {8.9, 10.8, 9.3},
  {10.6, 11.4, 9.1},
  {13.8, 12.4, 9.3},
  {15.1, 14.8, 9.8},
  {16.5, 16.5, 11.8},
  {18, 16.6, 15.7},
  {18.4, 17.8, 18.7},
  {18.2, 18.6, 21.2},
  {17.3, 19, 21.2},
  {15.8, 16.6, 18.4},
  {13.7, 14.1, 15.9},
  {12.4, 13.2, 13.9},
  {11.6, 12.5, 12.3},
  {11.7, 12.4, 11.2},
  {11.5, 12.2, 10.6},
  {11.2, 12, 9.9},
  {11.3, 11.9, 9.4},
  {11.3, 11.9, 9},
  {11.1, 11.6, 8.6},
  {11.2, 12.1, 8.6},
  {11.5, 11.7, 9.1},
  {11.2, 11, 9.1},
  {11.2, 11.3, 9.1},
  {11.5, 10.7, 9},
  {12.2, 10.6, 8.8},
  {14.2, 11, 8.8},
  {18.6, 12, 9.2},
  {19.1, 13.8, 10.5},
  {19.5, 16.3, 12.6},
  {19.4, 18.7, 15.9},
  {20.5, 19.3, 18.8},
  {20.1, 20, 21.3},
  {18.7, 19.4, 21.7},
  {16, 17.6, 18.8},
  {14.6, 15.3, 16.4},
  {14, 14.4, 14},
  {12.8, 13.5, 12.5},
  {12.7, 13.4, 11.5},
  {12.1, 13.7, 10.8},
  {11.5, 13.3, 10},
  {11.7, 12.5, 9.4},
  {11.4, 12.1, 8.8},
  {11.1, 11.6, 8.5},
  {10.5, 11.2, 7.8},
  {10.9, 11, 7.6},
  {10.8, 10.8, 7.1},
  {10.4, 10.8, 6.9},
  {10.4, 10.6, 6.5},
  {10.5, 10.8, 6.2},
  {13.7, 11.8, 6.6},
  {16.5, 14, 8.3},
  {17.6, 15.3, 11.3},
  {18.6, 16.9, 15.3},
  {18.2, 19.5, 18.8},
  {19.4, 20.1, 19.6},
  {19.9, 20.5, 21.5},
  {18.4, 20, 20.1},
  {15, 18, 18.3},
  {14.3, 16.3, 15.7},
  {13.3, 15.7, 13.5},
  {12.8, 15, 11.8},
  {12.1, 15.3, 10.5},
  {11.6, 15.8, 9.7},
  {12.1, 15.7, 8.9},
  {11, 14.7, 8},
  {11.4, 14.4, 7.4},
  {11.7, 14.1, 6.7},
  {11, 13.8, 6.2},
  {11, 13.9, 5.6},
  {10.9, 12.7, 5},
  {9.9, 12.4, 4.5},
  {8.2, 12.2, 3.9},
  {8.6, 11.6, 3.7},
  {11.8, 11.6, 3.9},
  {14.8, 12, 5},
  {15.8, 15.1, 8.8},
  {16, 17, 13},
  {15.9, 17.9, 16.6},
  {14.6, 18.3, 18.5},
  {13.1, 17.5, 17.6},
  {12.7, 15.8, 16.6},
  {11.5, 14.2, 15.1},
  {10.7, 13, 13.8},
  {10.2, 12.1, 10.7},
  {10.4, 11.2, 9.2},
  {10.2, 11.3, 7.9},
  {9, 10.2, 7.5},
  {7.7, 9.3, 6.9},
  {7, 8.9, 7},
  {7.2, 8.2, 7.4},
  {5.7, 7.9, 7.7},
  {5.4, 8.2, 7.7},
  {4.8, 7.9, 7.9},
  {4.9, 7.3, 7.1},
  {5.3, 7, 6.1},
  {4.4, 7, 5.4},
  {5.2, 7.6, 5.2},
  {7.4, 8.4, 5.2},
  {10.7, 9.1, 5.9},
  {11.3, 11.2, 8.6},
  {11.5, 11.8, 11.6},
  {11.8, 12.6, 13.4},
  {11.8, 13.2, 14.8},
  {12.5, 13.6, 15.6},
  {11, 12.8, 15.7},
  {9.6, 11.6, 14},
  {8.9, 10.5, 12.6},
  {8.6, 10.1, 10.8},
  {8.3, 9.8, 9.6},
  {7.9, 9.7, 9},
  {6.7, 9.7, 8.4},
  {6.9, 9.2, 7.6},
  {6.6, 9, 7.6},
  {6, 7.9, 7.2},
  {5.6, 7.5, 6.7},
  {5.2, 7.1, 6},
  {4.6, 6.6, 5.4},
  {4.6, 6.2, 4.6},
  {4.6, 6.1, 4.3},
  {4.4, 5.9, 3.8},
  {4.3, 5.7, 3.4},
  {6.4, 6.5, 3.5},
  {9.7, 6.7, 4.7},
  {10.8, 8.7, 6.8},
  {12.2, 10.9, 9.8},
  {13.1, 13.1, 13.2},
  {13.2, 14.6, 16},
  {13.6, 15.4, 17.1},
  {12.7, 14.9, 16.9},
  {11.1, 13.3, 13.8},
  {9.5, 11.4, 11.6},
  {8.2, 10.1, 10.7},
  {7.5, 9, 12.7},
  {6.4, 7.6, 11.8},
  {6.4, 6.9, 11.1},
  {5.6, 5.9, 10.3},
  {5.1, 5.4, 9.1},
  {4.5, 5.3, 8.1},
  {3.8, 5, 5.7},
  {3.5, 4.6, 4},
  {3, 4.1, 2.4},
  {1.3, 3.9, 1.3},
  {1, 4, 0},
  {0.9, 3.8, -0.7},
  {1, 3.5, -1.1},
  {1.9, 3.7, -0.9},
  {4.5, 4.3, 0.1},
  {5, 5.2, 4.7},
  {5, 5.7, 8.1},
  {5, 5.9, 8.2},
  {5.4, 6, 8.2},
  {5, 6.1, 8.4},
  {4.1, 5.8, 8.3},
  {2.6, 4.1, 7.6},
  {0.6, 2.9, 5.7},
  {-0.4, 2.6, 3.8},
  {-1.5, 2.1, 1.2},
  {-1, 1.4, -0.8},
  {-2.4, 0.6, -1.8},
  {-2.3, -0.1, -2.4},
  {-2.7, -0.5, -2.8},
  {-3, -0.6, -3.2},
  {-2.9, -0.7, -3.4},
  {-3.1, -1, -3.9},
  {-3.3, -1.4, -4.1},
  {-3.4, -1.6, -4.4},
  {-3.7, -1.7, -4.8},
  {-2.9, -1.6, -5},
  {-2.5, -1.4, -5.1},
  {-0.1, -0.9, -5},
  {3.5, -0.7, -4},
  {5, 2.4, -0.3},
  {5.5, 6, 3.4},
  {6.3, 7.4, 6.9},
  {7, 7.7, 9.9},
  {6.9, 8.1, 10.5},
  {6.2, 7.8, 10.4},
  {3.4, 5.8, 7.4},
  {1.4, 4.4, 4.9},
  {1.1, 3.7, 3.2},
  {0.1, 3.1, 2.4},
  {-0.3, 1.8, 1.5},
  {-0.1, 1.4, -0.2},
  {-0.2, 1.3, -1.5},
  {-1, 0.6, -2.2},
  {-0.9, 0.1, -2.8},
  {-2.3, 0.1, -3.3},
  {-2.7, 0, -3.5},
  {-2.8, -0.6, -4},
  {-3.7, -0.9, -4.5},
  {-4, -1.6, -4.6},
  {-3.8, -1.4, -4.8},
  {-3.6, -1.6, -5.1},
  {-1.8, -1.4, -5},
  {2.8, -0.6, -3.8},
  {4.6, 2.6, -0.4},
  {5.8, 5.6, 3.7},
  {6.5, 6.8, 6.9},
  {6.9, 8, 9.5},
  {7.2, 8.5, 10.9},
  {6.3, 8.4, 9.8},
  {4.4, 5.5, 7.6},
  {2.3, 3.7, 5.3},
  {1.8, 2.6, 2.8},
  {1.6, 1.9, 1.3},
  {0.6, 1.6, 0.2},
  {0.1, 1.1, -0.6},
  {0.4, 0.8, -1.6},
  {0.2, 0.7, -2.1},
  {-0.6, 0.8, -2.4},
  {-0.4, 0.3, -2.7},
  {-0.5, 0.4, -3.1},
  {-0.7, 0.4, -3.4},
  {-0.7, 0.3, -3.6},
  {-0.8, 0.5, -3.7},
  {-0.3, 0.7, -4},
  {0.2, 0.4, -4},
  {2.9, 0.9, -3.7},
  {6.1, 1.6, -1.9},
  {7.8, 4.4, 1.5},
  {8.9, 6.5, 4.7},
  {9.1, 8.2, 8.1},
  {9.8, 9.1, 10.4},
  {9.6, 10.2, 11.9},
  {10, 9.6, 12.8},
  {6.9, 7.4, 8.7},
  {5.9, 6.2, 5.8},
  {6.2, 6.5, 4.4},
  {5.9, 6.7, 3.6},
  {6.2, 6.1, 2.4},
  {5.5, 6, 1.2},
  {4.7, 5.8, 0.6},
  {5, 5.7, 0.4},
  {5.1, 5.5, -0.2},
  {4.9, 5.6, -0.3},
  {4.6, 5.2, -0.8},
  {5.2, 5, -1},
  {5.1, 5.1, -0.9},
  {5, 5.3, -1.1},
  {4.7, 4.8, -1.4},
  {5.7, 5.8, -1.6},
  {7.6, 7.2, -1.1},
  {9.9, 7.2, 0.3},
  {11.6, 8.6, 2},
  {12.2, 10, 4.8},
  {12.7, 10.3, 6.9},
  {13.1, 11, 8.5},
  {12.5, 10.1, 8.9},
  {10.6, 10.2, 8.4},
  {9.6, 10.1, 7.4},
  {8.7, 9.5, 5.5},
  {8.9, 9.8, 4.4},
  {8.1, 8.2, 3.6},
  {7.9, 8.6, 3.1},
  {7, 9, 1.9},
  {7.6, 8.6, 1.6},
  {6.9, 8, 1},
  {6.6, 8.1, 0.6},
  {6.7, 7.8, -0.1},
  {6.7, 8.2, -0.7},
  {5.7, 7.8, -1},
  {5.5, 7.2, -1.3},
  {5.8, 6.8, -1.6},
  {4.6, 6.2, -1.9},
  {5, 6, -1.9},
  {7, 6.5, -1.8},
  {11.4, 7.3, -0.9},
  {13, 10.7, 2.2},
  {13.6, 11.6, 8.5},
  {14.4, 13.9, 12.6},
  {14.9, 14.9, 15.3},
  {14.5, 14.5, 17.6},
  {12.8, 13.9, 16.9},
  {10, 10.7, 12.2},
  {7, 8.6, 8.1},
  {6.3, 7.5, 5.4},
  {5.4, 7, 3.8},
  {5.8, 6.6, 2.5},
  {5.4, 6.1, 1.7},
  {4.6, 5.7, 1.2},
  {4.2, 5.3, 0.6},
  {3.6, 4.9, 0.3},
  {4.3, 4.7, -0.5},
  {3.5, 4.1, -0.5},
  {2.9, 4.5, -1.1},
  {3, 3.9, -1.2},
  {3.3, 3.4, -1.7},
  {3.9, 3.1, -1.7},
  {3.9, 3.2, -1.7},
  {5.7, 3.3, -1.7},
  {8.7, 4.2, -0.8},
  {10.3, 6.9, 2.8},
  {11.9, 9.8, 7.2},
  {12.3, 11.7, 10.8},
  {11.5, 12.7, 13.9},
  {11.3, 12.8, 15.2},
  {10.5, 12.5, 14.2},
  {8.5, 10.2, 11.6},
  {8.1, 8.8, 8.2},
  {8.9, 8.5, 6.8},
  {8.3, 8.2, 6.2},
  {8.1, 7.2, 5.2},
  {7.2, 6.6, 4},
  {7.2, 6.3, 2.9},
  {7.4, 6.2, 2.1},
  {6.9, 5.9, 1.9},
  {6.3, 5.5, 1.4},
  {5.9, 5.5, 1.2},
  {5.5, 5.3, 0.7},
  {5.7, 5, 0.2},
  {4.6, 4.7, 0.5},
  {4.2, 4.3, 0.1},
  {4, 4.4, 0.5},
  {5.8, 4.4, 0.9},
  {10.2, 5.4, 1.4},
  {11.8, 7.1, 3.8},
  {11.9, 9.6, 5.8},
  {13.4, 9.6, 9.3},
  {13.3, 10.7, 13.2},
  {12.8, 10.8, 14.9},
  {11.8, 12, 15.8},
  {10.3, 9.5, 12.6},
  {8.3, 8.5, 9.7},
  {7.2, 8.5, 7.5},
  {7.3, 8.2, 5.9},
  {6.5, 7.3, 4.8},
  {6.7, 7, 4.3},
  {6.4, 6.9, 3.5},
  {5.4, 6.9, 2.8},
  {5.4, 7.3, 2.1},
  {5.5, 6.4, 1.4},
  {5.4, 7.7, 0.6},
  {5.7, 7, 0.1},
  {5.9, 7.8, 0.1},
  {5.8, 8.3, -0.3},
  {6.7, 7.3, -0.5},
  {7, 6.9, -0.4},
  {8, 6.1, -0.1},
  {10.7, 7.8, -0.2},
  {11.1, 9.5, 2.7},
  {12.2, 12, 6.3},
  {13, 13.1, 11.1},
  {12.7, 14.7, 16},
  {12.7, 14.7, 16.5},
  {10.9, 14.4, 15.9},
  {8, 11.1, 12.3},
  {7.2, 9.9, 10.8},
  {7.1, 8.8, 6.9},
  {6.3, 7.9, 5.4},
  {6.3, 7.2, 5.2},
  {5.5, 6.6, 4.6},
  {5.5, 6.2, 4.4},
  {6, 5.3, 4.9},
  {5.9, 4.9, 5.4},
  {5.3, 4.7, 5.4},
  {4.8, 4.7, 5.3},
  {4, 4.6, 5.2},
  {3.7, 4.4, 4.8},
  {3.3, 4.1, 3.5},
  {2.2, 3.7, 2.7},
  {2.1, 3.9, 2},
  {3.8, 4.3, 2.1},
  {5.2, 4.5, 3.3},
  {6, 5.1, 5.1},
  {6.2, 5.4, 6.7},
  {6.2, 5.7, 7.6},
  {6.3, 6.3, 8.1},
  {5.7, 5.7, 8.3},
  {5, 5.6, 7.8},
  {4.2, 5.4, 7.1},
  {3.3, 4.7, 6.1},
  {2.9, 4.7, 4.6},
  {2.7, 4.1, 4},
  {2.2, 3.8, 3.1},
  {1.8, 3.1, 2.1},
  {1.7, 2.9, 1.1},
  {1.4, 2.7, 0.6},
  {1.3, 2.4, -0.2},
  {1.6, 2, -0.4},
  {2.9, 1.5, -0.8},
  {3.5, 1.4, -0.9},
  {3.2, 1.3, -1.1},
  {3.1, 1.1, -0.9},
  {2.4, 1.7, -0.8},
  {2.8, 2.2, -0.9},
  {2.9, 1.9, -0.5},
  {5.8, 2.1, -0.1},
  {7.1, 3.9, 2.2},
  {8.6, 6.2, 5.8},
  {9.9, 7.1, 8.8},
  {10.2, 9.3, 11.8},
  {10.4, 9.3, 13.3},
  {8.2, 8.8, 13},
  {6.9, 8.8, 9.7},
  {5.8, 8.8, 6.8},
  {6.7, 9.5, 4.8},
  {5.4, 8.8, 3.8},
  {6.3, 8.6, 2.6},
  {5.4, 9.1, 2.3},
  {4.9, 8.6, 1.3},
  {4, 7, 0.8},
  {2.9, 6.8, 0.5},
  {2.7, 6, 0},
  {1.6, 5.2, -0.7},
  {1.3, 4.5, -1.1},
  {0.9, 4.4, -1.6},
  {0.9, 3.7, -2.2},
  {0.7, 4.1, -2.2},
  {1, 3.1, -2.6},
  {2.3, 3.3, -2.4},
  {7.5, 4, -2},
  {9.5, 5.9, 1.7},
  {10.3, 9.1, 5.7},
  {10.7, 10.6, 9.7},
  {11.2, 11.9, 12.3},
  {11, 12, 13.8},
  {9.8, 11.3, 12.9},
  {7.2, 9.9, 10.6},
  {4.6, 7.9, 7.6},
  {4.2, 6.9, 5.3},
  {3.5, 5.9, 3.3},
  {2.7, 4.9, 2.1},
  {2.5, 4.4, 1.3},
  {2.2, 3.9, 0.4},
  {2.3, 3.7, 0},
  {1.7, 3.8, -0.5},
  {2.2, 3.4, -0.8},
  {2.3, 3.2, -1},
  {3.4, 3.6, -1.2},
  {3.6, 3.6, -0.8},
  {3.6, 3.7, -0.5},
  {2.8, 3.4, -0.6},
  {3.5, 3.1, -1.1},
  {4.5, 3.6, -1.1},
  {9, 4.5, -0.8},
  {10.6, 6.5, 2.3},
  {11.6, 9.4, 6.9},
  {11.6, 10.6, 11},
  {11.4, 11.4, 13.8},
  {10.4, 12.1, 14.9},
  {9.9, 11.3, 13.6},
  {8.4, 8.7, 10.6},
  {6.8, 7.7, 7.2},
  {6.8, 7.1, 5.3},
  {6, 6.4, 3.7},
  {6.7, 6, 3},
  {6.8, 5.6, 1.9},
  {6, 5.1, 1.5},
  {6.6, 4.8, 1},
  {5.9, 4.9, 0.8},
  {5.1, 5.3, 0.6},
  {4.3, 5.8, 0.5},
  {4.9, 5.9, 0.5},
  {4.5, 5.7, -0.1},
  {3.9, 5.6, 0},
  {3.5, 5.3, 0.1},
  {3.4, 5.2, 0},
  {5, 4.8, -0.2},
  {7.5, 5.4, 0.6},
  {8.6, 6.5, 3.9},
  {9.5, 8.6, 6.2},
  {10.4, 9.7, 10.4},
  {10.3, 10.9, 12.5},
  {10.3, 11.7, 13.5},
  {9.8, 10.9, 12.9},
  {7.4, 8.6, 10.8},
  {5.6, 7.2, 8.1},
  {5.6, 6.6, 6.2},
  {6, 6.2, 4.6},
  {5.5, 5.9, 3.3},
  {5.3, 6.6, 2.3},
  {5.5, 6.9, 2.2},
  {6.4, 6.3, 1.6},
  {6.3, 5.9, 1.5},
  {6.3, 5.9, 2.1},
  {6.1, 5.7, 1.8},
  {5.6, 5.7, 1.6},
  {6.5, 5.8, 2.1},
  {6.5, 5.9, 2.7},
  {6.4, 6, 3.2},
  {7, 6.2, 3.6},
  {7.6, 6.4, 4},
  {8.5, 6.6, 4.6},
  {9.2, 7, 5.8},
  {8.3, 7.9, 7.2},
  {9.3, 8.7, 8.9},
  {10, 9.6, 10.2},
  {10, 10.1, 13.2},
  {9.2, 9.8, 13.1},
  {9.1, 10, 11.8},
  {8.7, 8.8, 10.5},
  {8.7, 8.7, 9.7},
  {8.7, 8.6, 9},
  {8.6, 8.5, 8.4},
  {8.6, 8.2, 8.1},
  {8.4, 8, 7.9},
  {8.3, 8.1, 7.5},
  {8.3, 8.1, 6.6},
  {8.2, 8, 6.5},
  {8.2, 7.7, 6.1},
  {7.9, 7.8, 6.4},
  {8, 7.7, 6.6},
  {7.6, 7.7, 6.6},
  {7.5, 7.7, 6.7},
  {8.5, 7.7, 6.2},
  {9.5, 7.9, 6.4},
  {10.3, 8.1, 6.8},
  {11.3, 8.6, 7.8},
  {11.9, 9.1, 8.9},
  {12, 10.2, 10.7},
  {12, 11.5, 12.1},
  {12.4, 12.7, 12.8},
  {12, 12.5, 13.5},
  {10, 11.7, 12.9},
  {8.2, 10.2, 10.4},
  {8.1, 9.2, 8.6},
  {7.6, 8.7, 7.4},
  {8.9, 8.7, 6.6},
  {9.2, 9.9, 6.9},
  {9, 9.3, 7.1},
  {9, 9, 7.3},
  {9.1, 8.8, 7.3},
  {9, 8.5, 7.4},
  {8.6, 8.2, 7.5},
  {8.5, 8.1, 7.5},
  {8.5, 8.2, 7.4},
  {8.7, 8.2, 7.6},
  {8.7, 8.2, 7.5},
  {8.8, 8.2, 7.5},
  {8.9, 8.4, 7.7},
  {9.1, 8.7, 7.9},
  {9.8, 9.1, 8.6},
  {10.7, 9.2, 9.4},
  {10.9, 9.8, 10.5},
  {10.8, 9.5, 11.4},
  {9.8, 10, 11.8},
  {9.3, 9.8, 12.1},
  {9, 9.8, 11.4},
  {8.9, 9.8, 10.8},
  {8.4, 9.6, 10.4},
  {7.8, 9.2, 10.2},
  {8, 9.4, 10},
  {7.3, 9.4, 9.8},
  {6.1, 9.4, 9.6},
  {5.9, 9.1, 9.4},
  {5.7, 9.1, 9.4},
  {5.2, 8.9, 9.1},
  {5.2, 9, 8.8},
  {5.1, 9, 8.1},
  {6.1, 8.8, 7.9},
  {5.1, 8.8, 7.8},
  {5, 8.8, 7.7},
  {4.8, 8.8, 7.5},
  {5.2, 8.7, 7.3},
  {8, 8.8, 7.3},
  {9.4, 9, 7.8},
  {10.5, 9.1, 8.3},
  {11.1, 9.6, 9.5},
  {11.7, 9.9, 10.5},
  {11.4, 10.8, 11.8},
  {10, 11.2, 12.5},
  {8.5, 8.7, 11.2},
  {7.2, 8.4, 10.2},
  {6.2, 7.8, 9},
  {5.7, 8.1, 8.6},
  {5.3, 7.7, 7.8},
  {6.3, 8, 7.5},
  {6.7, 8.2, 7.4},
  {6.9, 7.8, 7.1},
  {6.6, 7.5, 7},
  {6.1, 6.8, 6.6},
  {6.4, 6.7, 6.8},
  {6.5, 7, 6.8},
  {6.3, 7.1, 6.9},
  {6.2, 7.1, 6.7},
  {6.2, 7, 6.8},
  {6.1, 6.9, 6.9},
  {6.2, 7.1, 7},
  {6.3, 7.1, 7.3},
  {6.6, 7.5, 7.7},
  {7.1, 8.1, 8.8},
  {7.5, 9, 9.9},
  {8.4, 10.3, 11},
  {9.6, 11.3, 13.3},
  {8.9, 10.1, 12.4},
  {6.5, 7.5, 9.9},
  {4.7, 6.1, 8.4},
  {4.3, 5.4, 7.3},
  {4.2, 5.5, 6.2},
  {4.8, 5.6, 6.3},
  {4.9, 6.1, 6.2},
  {4.7, 6.2, 5.5},
  {5, 5.8, 5.4},
  {5.1, 5.7, 5.6},
  {5, 5.6, 5.6},
  {5, 5.6, 5.7},
  {5.2, 5.5, 5.7},
  {5.2, 5.4, 5.8},
  {5.1, 5.1, 5.8},
  {4.9, 5.1, 5.6},
  {4.7, 5.1, 5.6},
  {5, 5.4, 5.4},
  {5.4, 5.3, 5.6},
  {5.6, 6, 6},
  {6.2, 6.7, 7.3},
  {8, 7.1, 10.1},
  {8.2, 7.7, 11.1},
  {6.5, 7.8, 10.7},
  {5.6, 7.6, 10.3},
  {5.2, 6.5, 9.4},
  {5.1, 6.3, 8.9},
  {5.1, 5.9, 8.2},
  {5.1, 5.7, 7.5},
  {4.9, 5.5, 7.3},
  {4.6, 5.5, 7},
  {4.3, 5.1, 6.9},
  {4.2, 4.8, 6.8},
  {4, 4.6, 6.7},
  {3.9, 4.5, 6.3},
  {3.7, 4.4, 6},
  {3.5, 4.1, 5.8},
  {3.3, 4, 5.6},
  {3.1, 4.3, 5.4},
  {2.9, 4.4, 5.2},
  {2.7, 4.2, 4.9},
  {2.9, 4.6, 4.8},
  {4.2, 5, 4.8},
  {6.3, 6, 5.6},
  {8.7, 7.5, 7.7},
  {9.6, 9.2, 10},
  {9.9, 10.6, 12},
  {9.7, 11, 12.6},
  {8.8, 10.4, 12},
  {6.6, 8.2, 9.1},
  {6, 7.4, 6.5},
  {5.4, 6.5, 4.9},
  {4.3, 5.3, 3.4},
  {4.4, 4.2, 2.5},
  {2.1, 3.7, 1.6},
  {0.7, 3.5, 1},
  {1.7, 3.1, 0.6},
  {1.7, 3, 0.5},
  {1.5, 3.1, 0.5},
  {1.3, 2.2, 0.3},
  {0.2, 2.2, 0.1},
  {0.5, 2.2, -0.4},
  {0.6, 1.6, -0.9},
  {1.1, 1, -1.1},
  {1.3, 0.9, -1.4},
  {0.9, 1.3, -1.4},
  {3.4, 2.7, -1},
  {5.4, 4.1, 0.4},
  {6.4, 5.6, 3.3},
  {6.1, 6.1, 6.2},
  {7.4, 6.8, 7.7},
  {7.2, 6.1, 8.8},
  {6.3, 5.9, 9},
  {3.9, 4.4, 7.6},
  {3, 3.2, 5},
  {2.6, 3, 3.2},
  {1.9, 2.9, 2.2},
  {2.4, 2.5, 1},
  {2.6, 2.3, 0.5},
  {3.3, 2.2, 0.1},
  {3.1, 2.4, -0.1},
  {3.9, 2.5, -0.4},
  {4, 2.8, -0.8},
  {3.9, 2.7, -0.7},
  {4.2, 2.8, -0.1},
  {4.1, 2.6, 0.2},
  {4.5, 2.9, 0.5},
  {4.3, 2.8, 0.4},
  {4.7, 2.9, 0.4},
  {5.3, 3.3, 0.9},
  {5.4, 3.4, 1.8},
  {6.1, 4.1, 3.3},
  {6.7, 5.2, 4.8},
  {7.3, 4.8, 7.2},
  {7.1, 6.2, 9.2},
  {6.5, 5.9, 10.1},
  {6.4, 6.2, 10},
  {5.6, 5.9, 9.4},
  {5.5, 5.1, 7.9},
  {6, 5.2, 6.9},
  {5.6, 4.5, 6.5},
  {5.7, 4.6, 6.3},
  {6.4, 4.4, 5.8},
  {6.6, 4.4, 5.5},
  {6.4, 4.6, 5.6},
  {6.6, 4.6, 5.7},
  {6.6, 4.5, 5.6},
  {6.1, 4.7, 5.5},
  {5.3, 4.5, 5.6},
  {5.7, 4.7, 5.6},
  {5.4, 4.9, 5.6},
  {5.5, 4.7, 5.3},
  {6.1, 4.9, 5.2},
  {6.7, 5.3, 5.2},
  {7.4, 5.6, 5.7},
  {8.1, 6.4, 6.5},
  {8.6, 6.7, 7.8},
  {9.4, 7, 9.4},
  {8.7, 8.2, 10.1},
  {9.1, 7.6, 10.5},
  {9.2, 7.8, 11},
  {9.5, 7.6, 10.8},
  {8.6, 7.5, 9.7},
  {8.2, 7.6, 8.7},
  {8.4, 7.7, 8},
  {8.7, 7.7, 7.5},
  {8.2, 8, 6.8},
  {7.5, 7.7, 5.9},
  {7.2, 7.5, 5},
  {6.6, 7.7, 4.3},
  {6.8, 7.6, 3.7},
  {6.3, 7.9, 3.4},
  {6.7, 7.5, 3.2},
  {5.8, 7.3, 2.8},
  {5.9, 7.1, 2.8},
  {5.9, 6.5, 3},
  {5.5, 6.6, 3.4},
  {6.2, 6.8, 3.8},
  {8.6, 7.3, 4.4},
  {10.4, 8.7, 4.8},
  {11.4, 9.8, 5.6},
  {12.3, 11, 8.3},
  {13.1, 12.3, 11.9},
  {12.9, 12.5, 14.8},
  {11.5, 11.9, 14.6},
  {8.7, 9.5, 11.1},
  {7.3, 8.4, 8.6},
  {6.9, 7.5, 7.8},
  {6.4, 7.2, 7.8},
  {6.1, 7.1, 7.3},
  {5.4, 6.7, 6.4},
  {5.6, 6.8, 5.9},
  {5.4, 6.5, 5.4},
  {4.7, 6.3, 5},
  {4.9, 5.8, 4.6},
  {4.8, 5.8, 4.3},
  {4.7, 5.7, 4},
  {4.1, 5.5, 3.6},
  {3.8, 4.8, 3.4},
  {4.1, 4.8, 3.2},
  {4.1, 4.6, 2.9},
  {4.8, 5, 2.9},
  {7.3, 5.6, 2.8},
  {9.2, 5.3, 3},
  {10, 7.9, 3.4},
  {9.9, 9.3, 4.7},
  {10.5, 10.1, 7.6},
  {10.1, 10.1, 11.2},
  {9.1, 9.6, 12.7},
  {5.7, 7.4, 9.2},
  {4.2, 6.1, 7.3},
  {3.6, 5.4, 5.4},
  {3.2, 4.9, 4.1},
  {2.5, 4.4, 3.4},
  {2.1, 4.4, 3.9},
  {2.5, 4.2, 4.6},
  {3, 4.2, 5.1},
  {3.6, 4.3, 5.2},
  {3, 4, 5.2},
  {3.4, 3.7, 5.1},
  {3.5, 3.4, 4.9},
  {2.9, 3.4, 4},
  {3.1, 3.1, 3.8},
  {2.6, 2.9, 3.5},
  {2.3, 2.2, 3.2},
  {3.2, 2.5, 2.9},
  {4.7, 2.9, 2.8},
  {6.2, 3.8, 2.9},
  {7.6, 4.8, 3.1},
  {7.4, 5.7, 3.7},
  {7.4, 6.4, 4.7},
  {7.6, 6.7, 7.1},
  {7.1, 7.1, 9},
  {4, 5.8, 7.3},
  {2.4, 4.5, 5.4},
  {2, 4, 3.9},
  {3.1, 3.3, 2.8},
  {2.8, 3, 2},
  {2.2, 2.8, 1},
  {2.2, 2.4, 1.4},
  {1.8, 2.2, 2.6},
  {1.3, 2, 2.8},
  {1, 2.1, 3},
  {1, 2.1, 3.1},
  {1.6, 1.9, 3.1},
  {1.5, 1.6, 3.1},
  {1.5, 1.6, 3},
  {1.8, 1.6, 2.8},
  {1.6, 1.4, 2.6},
  {2.2, 0.4, 2},
  {5.8, 2.4, 1.7},
  {8.3, 2.3, 1.6},
  {9.4, 4.4, 2},
  {9.9, 5.9, 3},
  {9.8, 7.5, 5.9},
  {9.3, 9, 9.1},
  {8.6, 8.3, 10.2},
  {5.1, 5.8, 6.4},
  {4.1, 4.9, 4.4},
  {4.9, 4.9, 2.9},
  {6.4, 5.3, 2},
  {6, 5.5, 1.1},
  {7, 5.6, 0.6},
  {7, 5.5, 0.2},
  {6.2, 5.4, -0.1},
  {6.6, 6.2, -0.4},
  {7.4, 5.8, -0.6},
  {7.3, 5.5, -1},
  {7.1, 4.8, -1},
  {6.9, 5.2, -1.2},
  {5.3, 4.7, -1.5},
  {5.2, 4.9, -1.7},
  {3.6, 4.4, -1.9},
  {3.9, 4.8, -1.8},
  {6.6, 5.6, -1.8},
  {9.2, 6.3, -0.1},
  {9.9, 7.8, 3.3},
  {10.4, 9.6, 6.7},
  {10.3, 10.4, 10.1},
  {10.3, 11, 13},
  {9.3, 10.5, 11.5},
  {6.5, 8, 7.1},
  {4.2, 6.4, 4.6},
  {3.6, 5.6, 3},
  {3.1, 4.8, 1.9},
  {2.8, 4.3, 1.1},
  {2.4, 4.5, 0.6},
  {2.5, 4.2, 0},
  {2.1, 3.9, 0},
  {2.5, 3.6, -0.8},
  {2.6, 3.3, -0.8},
  {3.1, 2.9, -1.2},
  {2.6, 2.8, -1.8},
  {1.9, 2.4, -1.7},
  {1.5, 2.1, -2.2},
  {1, 1.8, -2.6},
  {0.7, 1.7, -2.6},
  {1.2, 1.5, -2.3},
  {3.5, 2.2, -2.1},
  {5.7, 3.4, -1.1},
  {7, 5.1, 1.6},
  {7.6, 6.6, 4.8},
  {7.4, 8.2, 8.1},
  {7.3, 8.4, 10.6},
  {7.1, 7.9, 9.7},
  {3.4, 5.5, 5.6},
  {2, 3.9, 3.2},
  {1.4, 3, 1.9},
  {0.9, 2.6, 0.6},
  {0.6, 2.2, 0},
  {0.4, 1.8, -0.4},
  {0.3, 1.8, -1},
  {0, 1.5, -1.5},
  {0, 1, -1.7},
  {-0.1, 0.8, -2.1},
  {-0.6, 0.6, -2.2},
  {-0.3, 0.3, -1.9},
  {-0.8, 0.2, -1.9},
  {-0.7, -0.1, -2.2},
  {-1.1, -0.5, -2.5},
  {-1.1, -0.6, -2.3},
  {-1.1, -0.6, -2.3},
  {1.2, -0.2, -2.3},
  {3.3, 0.8, -1.9},
  {4.5, 4.1, -0.7},
  {4.9, 5.7, 1.7},
  {5.2, 6, 4.7},
  {5.2, 6.5, 7.1},
  {4.3, 5.4, 7.6},
  {2.8, 3.4, 4.3},
  {2.6, 2.2, 2.1},
  {2.6, 1.7, 0.5},
  {2.6, 2.4, 0.1},
  {2.6, 2.5, -0.5},
  {2.4, 2.6, 0.1},
  {2.2, 2.3, 0.5},
  {1.6, 2.2, 0.8},
  {0.7, 1.9, 0.9},
  {0.4, 1.9, 0.7},
  {0.6, 1.3, -0.1},
  {-0.1, 0.9, -0.8},
  {-0.5, 0.8, -1.2},
  {-0.3, 0.8, -1.4},
  {0.1, 1.2, -1.2},
  {0.7, 1.8, -1},
  {1.3, 2.2, -0.9},
  {1.6, 2.6, -0.7},
  {2.9, 1.1, 0.3},
  {4.9, 1.6, 2.2},
  {5.5, 2.4, 4},
  {7.7, 2.6, 6.2},
  {6.8, 3, 6.7},
  {5.6, 3.1, 6.5},
  {5.1, 2.9, 6.3},
  {4.9, 3, 5},
  {5, 3, 4.3},
  {5.5, 2.9, 4.2},
  {5.7, 3.1, 3.9},
  {5.7, 2.6, 3.9},
  {5.4, 2.8, 3.8},
  {5.1, 2.5, 3.7},
  {5.2, 2.8, 3.7},
  {4.8, 2.8, 3.6},
  {4.4, 2.8, 3.6},
  {4.7, 3, 3.6},
  {4.8, 2.8, 3.5},
  {4, 3, 3.5},
  {3.6, 3.1, 3.1},
  {3.8, 3, 3.1},
  {3.5, 2.9, 3.2},
  {3.8, 3, 3.6},
  {5, 3.6, 4.2},
  {5.9, 3.9, 5.2},
  {5.2, 4.8, 6.3},
  {4.6, 5.6, 7.9},
  {5.3, 5.1, 8.9},
  {4.7, 5.2, 8.2},
  {3.8, 4.6, 6.8},
  {3.3, 4.7, 5.1},
  {2.9, 4, 4.4},
  {2, 3.3, 2.9},
  {2, 3.2, 2},
  {1.9, 2.9, 1.3},
  {2, 2.9, 1.2},
  {2.4, 2.7, 0.8},
  {2.2, 2.7, 0.4},
  {2.3, 2.7, 0.4},
  {2.1, 3.6, 0.8},
  {2.6, 3.3, 1.4},
  {2.9, 2.8, 1.8},
  {3.5, 3.5, 2.3},
  {3.5, 4.3, 2.5},
  {3.1, 3.9, 2.4},
  {3.7, 5, 2.2},
  {5, 5, 2.1},
  {6.2, 5.1, 2.2},
  {7, 5.8, 2.8},
  {7, 7, 4.4},
  {8.4, 7.7, 6.3},
  {7.8, 7.9, 9},
  {7.9, 7.7, 9.4},
  {5.2, 6, 7.2},
  {3.7, 5.4, 5.1},
  {4, 4.7, 3.9},
  {4.3, 5.2, 4.4},
  {4.5, 5.3, 4.7},
  {4.5, 5.2, 4.5},
  {4.8, 5, 4.6},
  {4.4, 5, 4.4},
  {5.3, 5, 4.6},
  {5.5, 4.7, 4.8},
  {5.8, 4.6, 4.6},
  {5.5, 4.8, 4.6},
  {5.9, 4.7, 4.6},
  {6.1, 4.3, 4.6},
  {6.4, 4.6, 4.6},
  {7.2, 4.5, 4.7},
  {7, 4.5, 4.7},
  {7.4, 4.7, 4.9},
  {8.1, 5, 5.2},
  {8.3, 5, 5.4},
  {8.1, 5.4, 5.7},
  {8.8, 5.8, 6},
  {8.9, 6.2, 6.3},
  {8.9, 5.9, 6.6},
  {9.1, 6, 6.5},
  {9.2, 6.3, 6.4},
  {8.8, 6.4, 6.2},
  {9.3, 6.6, 6.1},
  {8.3, 6.7, 6.2},
  {8.1, 6.9, 6.2},
  {7.6, 6.8, 6.4},
  {6.7, 6.8, 6.3},
  {6.7, 7.5, 5.9},
  {6.8, 7, 6},
  {7.3, 6.6, 6.1},
  {7.4, 7, 6.3},
  {7.2, 7, 6.4},
  {7.2, 6.7, 6.4},
  {7.4, 7, 6.4},
  {7.2, 7.2, 6.5},
  {7.4, 7.1, 6.5},
  {7.9, 7.3, 6.7},
  {8, 7.6, 6.9},
  {8.1, 7.9, 7.5},
  {7.9, 7.8, 8.1},
  {7.7, 7.9, 8.6},
  {7.8, 8.4, 9.2},
  {8.1, 8.5, 9.6},
  {7.8, 8.3, 9.5},
  {7.6, 8.2, 9.1},
  {7.5, 8.3, 8.8},
  {7.5, 8.2, 8.5},
  {7.4, 8.2, 8.4},
  {7.4, 8.2, 8.4},
  {7.5, 8.2, 8.2},
  {7.5, 8.2, 8.2},
  {7.2, 8.6, 7.9},
  {7.1, 8.3, 7.8},
  {7.1, 8.2, 7.7},
  {7.4, 8.2, 7.6},
  {7.7, 8.1, 7.4},
  {7.7, 8.1, 7.3},
  {7.5, 8.3, 7.3},
  {7.6, 8.2, 7.5},
  {7.8, 8.3, 7.3},
  {8, 8.4, 7.4},
  {8.1, 8.4, 7.7},
  {8.2, 8.4, 8.1},
  {8.2, 8.3, 8.4},
  {8.4, 8.3, 9},
  {9.4, 8.7, 9.1},
  {8.5, 8.5, 9.3},
  {8.2, 8, 8.8},
  {8.1, 7.8, 8},
  {8, 7.5, 7.7},
  {8.1, 7.3, 7.5},
  {7.7, 6.9, 7.2},
  {7.8, 7.2, 7},
  {7.2, 7, 6.7},
  {7.2, 6.8, 6.5},
  {6.8, 6.8, 6.5},
  {6.2, 6.6, 6.1},
  {5.7, 6.2, 5.7},
  {5.1, 5.7, 5.1},
  {4.6, 5, 4.2},
  {4.8, 3.5, 3.7},
  {4.9, 3.3, 3.5},
  {4.7, 3.1, 3.4},
  {4.5, 3.5, 3.3},
  {4.5, 3.3, 3.4},
  {4, 3.2, 3.5},
  {5.1, 3.5, 3.8},
  {6.3, 4.1, 4.8},
  {5.9, 4.3, 6.2},
  {5.9, 4.7, 7.8},
  {5.8, 4.7, 7.9},
  {3.8, 4.4, 7.1},
  {2.3, 4.1, 6.5},
  {2.5, 3.7, 6.1},
  {2.3, 2.7, 5.9},
  {2.1, 2.7, 5.9},
  {1.4, 3, 5.5},
  {1.3, 3, 5},
  {1.6, 3, 4.6},
  {1.1, 2.7, 4.1},
  {0.9, 2.6, 3.5},
  {1.1, 2.2, 3.1},
  {1.3, 2.2, 3.1},
  {1, 2.1, 3.1},
  {0.7, 1.9, 3},
  {1, 2, 3},
  {1.1, 1.8, 2.8},
  {1.2, 2.1, 2.7},
  {3.1, 3.4, 3.2},
  {4.1, 4.3, 3.7},
  {5.4, 5.9, 4.4},
  {5.2, 7.1, 5.2},
  {6.2, 7.1, 6.5},
  {6.3, 6.5, 7.9},
  {5.8, 4.2, 8.8},
  {2.2, 3, 5.7},
  {1.1, 2.2, 4.1},
  {0.3, 1.7, 2.8},
  {0, 1.8, 1.6},
  {-0.4, 1.3, 0.7},
  {-0.4, 0.9, 0.2},
  {-0.7, 0.3, -0.2},
  {-0.9, 0, -0.6},
  {-1.3, -0.3, -0.8},
  {-1.5, -0.6, -1},
  {-1.7, -0.7, -0.9},
  {-1.6, -0.8, -0.6},
  {-2.2, -0.9, -1},
  {-2.4, -1.2, -1.4},
  {-2.7, -1.4, -1.8},
  {-2.9, -1.5, -1.9},
  {-2.6, -1.5, -2.1},
  {-0.9, -1.3, -2.4},
  {1.3, -0.4, -2.4},
  {1.7, 1.1, -2},
  {3, 2.1, -0.3},
  {3.1, 3, 2.2},
  {3.6, 3.9, 4.8},
  {3.5, 2.7, 4.6},
  {0, 0.8, 1.7},
  {-0.9, 0.1, 0.3},
  {-1.3, 0, -0.2},
  {-1.2, -0.2, -0.6},
  {-2, -0.2, -0.9},
  {-2, -0.5, -1.4},
  {-2, -0.4, -1.8},
  {-2.1, -1, -2},
  {-2.3, -0.8, -2.2},
  {-1.6, -1, -2.5},
  {-2.6, -1.1, -2.9},
  {-2.7, -1.2, -3.1},
  {-2.8, -1, -3.1},
  {-2.4, -1.5, -2.9},
  {-2.5, -1.2, -3.3},
  {-2.1, -0.4, -3.2},
  {-0.7, -0.1, -2.6},
  {0.3, 0.7, -1.9},
  {1.8, 0.7, -1.1},
  {1.9, 2.2, 0.1},
  {2.2, 2.6, 2},
  {4.2, 3.2, 3.9},
  {5.4, 4.1, 5.8},
  {3.8, 3.1, 6},
  {1, 1.9, 2.9},
  {0.8, 1.4, 1.6},
  {0.4, 1.2, 0.5},
  {-0.3, 1.1, -0.1},
  {-0.1, 0.6, -0.5},
  {-0.6, 0.3, -0.9},
  {-0.3, 0.5, -1.4},
  {0, 0.4, -1.5},
  {0.1, 0.3, -1.8},
  {0, 0, -2},
  {-0.1, 0, -2.4},
  {-0.3, 0, -2.7},
  {-1, 0.3, -2.8},
  {-0.6, -0.1, -3.1},
  {-0.3, 0, -3.2},
  {-0.3, -0.1, -3.5},
  {0, 0.3, -3.4},
  {1.7, 0.3, -3.3},
  {4.2, 0.9, -2.3},
  {5.3, 4.2, 0.4},
  {7.1, 4.1, 3.1},
  {8.1, 6, 5.7},
  {8, 6.9, 7.5},
  {7.5, 5.8, 7.4},
  {2.6, 4, 2.9},
  {2, 3.5, 1.2},
  {1.8, 2.8, 0.2},
  {1.7, 2.8, -0.4},
  {1.6, 2.8, -0.8},
  {2.1, 2.1, -1.2},
  {1.9, 2, -1.5},
  {1.5, 2, -1.9},
  {1.5, 1.9, -2.1},
  {1.8, 1.3, -2.6},
  {1.2, 1.1, -2.7},
  {0.6, 1, -3},
  {0.3, 1, -3.3},
  {0.8, 0.9, -3.5},
  {0.8, 1.1, -3.6},
  {1, 0.7, -3.9},
  {1, 0.7, -3.8},
  {3.2, 1.9, -3.8},
  {6.1, 3.4, -2.7},
  {8.2, 5.5, 0.2},
  {9.2, 6, 3.3},
  {10.3, 6.2, 6},
  {11, 6.8, 7.9},
  {10, 6.9, 7.4},
  {4.7, 5.1, 3},
  {3.1, 4.2, 1.3},
  {3.1, 4, 0.3},
  {3.3, 3.2, -0.3},
  {3.2, 3.3, -0.8},
  {2.8, 2.9, -1.3},
  {2.2, 2.4, -1.5},
  {2.3, 2.7, -2},
  {2.3, 2.2, -2.4},
  {2.1, 2.1, -2.4},
  {2.5, 1.9, -2.8},
  {2.4, 1.7, -3},
  {2.6, 1.8, -3.1},
  {1.6, 1.2, -3.4},
  {1, 1.2, -3.5},
  {1.5, 0.7, -3.9},
  {1.8, 0.9, -3.9},
  {4.9, 1.2, -3.8},
  {7.7, 1.7, -2.3},
  {9.5, 4.8, -0.1},
  {9.6, 5.6, 2.4},
  {9.8, 6.4, 5.1},
  {9.4, 6.2, 7.5},
  {8.2, 5.4, 6.8},
  {5, 4.2, 3.3},
  {4.1, 3.4, 1.6},
  {3.8, 3, 0.5},
  {3.6, 2.9, 0},
  {2.8, 3.2, -0.5},
  {2.5, 3.1, -1.1},
  {2.4, 3, -1.3},
  {2.9, 2.6, -1.6},
  {2.1, 2.3, -1.9},
  {2, 2.2, -2.3},
  {2.3, 1.7, -2.4},
  {2.4, 1.6, -2.8},
  {2.3, 1.7, -3},
  {2.2, 1.8, -3.2},
  {2, 1.6, -3.3},
  {1.4, 1, -3.4},
  {2.4, 1, -3.7},
  {4.7, 1.6, -2.9},
  {7, 1.2, -2.1},
  {7.8, 4.3, 0.3},
  {6.7, 4.6, 1.4},
  {7, 4.3, 2.6},
  {6, 4.5, 3.7},
  {6, 4.7, 3.7},
  {4.8, 4, 3},
  {4.4, 3.9, 2.5},
  {4.4, 3.6, 1.9},
  {4.7, 3.5, 1.7},
  {4.4, 3.1, 1.6},
  {4, 2.8, 1.4},
  {3.7, 2.8, 1.2},
  {3.2, 2.7, 1},
  {3.1, 2.2, 1},
  {3.3, 2.6, 1.3},
  {2.8, 2.7, 1.5},
  {2.8, 2.7, 1.5},
  {2.6, 2.2, 1.7},
  {2.8, 2.6, 1.7},
  {2.8, 2.4, 1.7},
  {3.2, 2.5, 1.7},
  {3.1, 2.9, 1.8},
  {3.5, 3.2, 2.1},
  {3.6, 2.7, 2.9},
  {4.2, 3.3, 4},
  {4.5, 3.8, 5.4},
  {4.9, 4.5, 6.9},
  {5.1, 4.9, 7.4},
  {4.9, 4.5, 7},
  {4.5, 4.6, 6.4},
  {4.5, 4.4, 5.1},
  {4.4, 4.4, 4.3},
  {4.2, 4.4, 4},
  {4.1, 4.3, 3.9},
  {3.7, 4, 3.7},
  {4, 4.1, 3.5},
  {4.4, 3.6, 3.3},
  {4.4, 3.7, 2.9},
  {4.3, 3.4, 2.8},
  {4.1, 3.1, 2.7},
  {4.2, 3.5, 2.5},
  {4.1, 3.8, 2.4},
  {3.8, 4.1, 2.2},
  {3.5, 4.4, 2},
  {3.3, 4.7, 1.8},
  {3.4, 4.7, 1.8},
  {3.5, 4.9, 2.2},
  {2.9, 5.7, 2.8},
  {2.3, 5.8, 3.4},
  {2.3, 5.7, 4.7},
  {2.5, 5.8, 5.9},
  {2.6, 5.7, 6.2},
  {2.4, 5.6, 6.1},
  {1.7, 5.5, 5.6},
  {1.5, 4.9, 4.9},
  {1.1, 4.9, 4.5},
  {1.3, 4.5, 3.9},
  {1.3, 4.4, 3.4},
  {1.2, 4.3, 3},
  {1.2, 4.1, 2.4},
  {1.2, 3.9, 2.2},
  {1.2, 3.6, 2},
  {1.1, 2.6, 1.6},
  {0.7, 2, 1.1},
  {0, 1.7, 0.3},
  {-0.8, 1.1, -0.2},
  {-1.2, 0.9, -0.6},
  {-1.5, 0.7, -1.3},
  {-1.5, 0.8, -1.7},
  {-0.4, 1.1, -1.3},
  {0.1, 2.1, -1.5},
  {0.6, 2.9, -0.9},
  {1.1, 3.3, -0.2},
  {1.4, 3.7, 0.8},
  {1.8, 4.4, 2.3},
  {1.7, 5, 3.3},
  {1.4, 4.9, 3.8},
  {0.8, 4.4, 3.7},
  {1, 3.6, 3.1},
  {1.2, 2.7, 2.1},
  {1.1, 2.6, 1.1},
  {0.5, 2.4, 0.7},
  {0.2, 1.8, 0.8},
  {-0.5, 1.3, 0.5},
  {-1.5, 1.2, -0.2},
  {-2.4, 0.7, -0.9},
  {-2.3, 0.3, -1.4},
  {-3, -0.3, -1.9},
  {-3.3, -0.3, -2.6},
  {-3.5, -0.8, -2.9},
  {-3.6, -0.9, -3.2},
  {-3.9, -1.1, -3.6},
  {-4.3, -1.4, -4},
  {-4.1, -1.4, -4.4},
  {-1.7, -1.2, -4.3},
  {0.6, -0.6, -3.6},
  {1.8, 1, -1},
  {3.1, 2.2, 1.8},
  {3.4, 2.8, 4.2},
  {3.5, 3.6, 5.9},
  {2.8, 3.2, 5.6},
  {-0.8, 1.1, 1.4},
  {-2.4, 0.2, -0.1},
  {-2.7, -0.4, -1.3},
  {-3.2, -0.5, -2.1},
  {-3.3, -0.8, -2.8},
  {-3.3, -1.1, -3.5},
  {-3.1, -1.1, -3.7},
  {-3.1, -1.3, -4.1},
  {-3.2, -1.6, -4.4},
  {-3.2, -2, -4.5},
  {-3, -1.7, -5},
  {-2.7, -1.4, -5},
  {-2.2, -2.2, -5.1},
  {-2.7, -2.3, -4.9},
  {-2.8, -2.2, -5.1},
  {-3, -2.2, -5.3},
  {-1.9, -2, -5.7},
  {0.7, -1.2, -5.9},
  {3.5, -0.7, -4.9},
  {4.4, 2.3, -1.5},
  {5.5, 3.7, 0.9},
  {4.5, 4.1, 3.1},
  {4, 4.4, 4.9},
  {3.9, 2.8, 4.7},
  {0.5, 0.9, 1.6},
  {0, 0.1, -0.1},
  {-0.3, -0.1, -1.3},
  {0.2, 0, -2},
  {0.4, -0.1, -2.7},
  {0, -0.5, -3.3},
  {-0.7, -0.6, -3.8},
  {-0.5, -0.8, -4},
  {-0.9, -1.1, -4.5},
  {-1.1, -0.6, -4.8},
  {-1.1, -0.9, -5.1},
  {-1.7, -1, -5.5},
  {-1.8, -1.9, -5.4},
  {-1.8, -1.3, -5.8},
  {-1.6, -1.8, -6.1},
  {-2.8, -2.2, -6.3},
  {-3, -1.7, -6.4},
  {-1.3, -0.9, -6.3},
  {1.6, -0.3, -5.3},
  {2.7, 1.9, -1.7},
  {2.7, 2.5, 0.7},
  {3.8, 3, 3.3},
  {4.3, 3.5, 5.4},
  {4.2, 3.2, 5},
  {-0.2, 1.5, 1},
  {-1.3, 0.7, -0.6},
  {-1.9, 0.5, -2},
  {-1.7, 0.1, -2.7},
  {-1.9, 0, -3.4},
  {-2.1, -0.3, -4.1},
  {-1.9, 0.1, -4.6},
  {-2.1, -0.9, -5.1},
  {-1.9, -1.2, -5.5},
  {-1.7, -1.4, -5.8},
  {-1.7, -0.4, -6},
  {-1.1, -0.4, -6.1},
  {-1.3, 0, -6.2},
  {-0.5, -0.5, -6.4},
  {0.1, -0.3, -6.4},
  {0.4, 0.2, -6.5},
  {1, 0.2, -6.5},
  {3.2, 1.5, -6.2},
  {6.3, 2.3, -5.4},
  {7.7, 4.9, -1.6},
  {8.9, 5.7, 1.5},
  {8.7, 5.2, 4.6},
  {9.9, 6.4, 6.8},
  {9.5, 5.7, 6.6},
  {7.3, 3.6, 2.4},
  {6.8, 2.9, 0.3},
  {6.5, 2.8, -0.7},
  {5.6, 3, -1.8},
  {5.7, 3, -2.3},
  {5.1, 2.8, -2.8},
  {4.9, 2.8, -3.2},
  {4.6, 2.6, -3.7},
  {5, 2.6, -4.1},
  {3.8, 2.7, -4.4},
  {4.5, 2.4, -4.8},
  {3, 2.1, -4.9},
  {3.1, 2.1, -5.1},
  {2.9, 1.9, -5.4},
  {2.9, 1.1, -5.6},
  {2.7, 1.1, -5.9},
  {1.7, 1.1, -6.2},
  {3.8, 1.2, -5.8},
  {6.2, 2.8, -4.4},
  {7.8, 6, 0.1},
  {8.8, 7.1, 2.6},
  {10.3, 8.1, 6},
  {11, 8.4, 8},
  {9.8, 6.8, 7.2},
  {4.7, 5.7, 2.8},
  {3.7, 4.6, 0.6},
  {3.7, 4.4, -0.4},
  {3.5, 4.3, -1.2},
  {3.6, 4, -1.8},
  {3.3, 3.6, -2.1},
  {3.2, 3.6, -2.7},
  {2.6, 3.9, -2.7},
  {3.2, 3, -3.2},
  {2.7, 3, -3.6},
  {2.7, 3.3, -3.8},
  {2.5, 3, -4.4},
  {2.9, 2.2, -4.3},
  {2.3, 2.6, -4.4},
  {2.3, 2.5, -4.7},
  {1.6, 2.2, -5.1},
  {2.5, 2.4, -4.8},
  {5, 2.7, -4.7},
  {8, 3.3, -3.8},
  {9.3, 5.9, -0.1},
  {10.8, 7.5, 3.3},
  {10.8, 7.6, 6.6},
  {11.5, 7.7, 9.5},
  {10.5, 7.6, 8.4},
  {5.1, 6, 3.7},
  {4, 5, 1.5},
  {2.9, 4.4, 0.2},
  {2.6, 4.5, -0.7},
  {2.2, 4.3, -1.4},
  {2, 3.8, -2},
  {1.4, 3.4, -2.5},
  {1.5, 3, -3.2},
  {1.1, 2.1, -3.6},
  {0.7, 2.1, -3.6},
  {0.3, 1.8, -4.1},
  {0.1, 1.2, -4.5},
  {0.2, 1.3, -4.9},
  {0.1, 1, -5.5},
  {0.4, 0.8, -5.4},
  {0, 1.1, -5.7},
  {0.3, 1.4, -5.9},
  {2.8, 1.5, -5.4},
  {5.4, 2.8, -4.6},
  {6.2, 5.5, 0},
  {5.6, 5.1, 2.7},
  {5.7, 5.9, 5.8},
  {5.7, 6.3, 7.7},
  {5.1, 5.3, 7.4},
  {1.2, 3, 3.3},
  {0.1, 1.8, 0.6},
  {0, 0.9, -0.8},
  {-0.9, 0.7, -1.9},
  {-0.7, 0.3, -2.6},
  {-0.7, 0.1, -3.5},
  {-1.4, 0.2, -3.7},
  {-1.1, -0.1, -4.3},
  {-1.6, 0, -4.9},
  {-1.5, -0.4, -5.1},
  {-1.4, -0.5, -5.3},
  {-1.3, -0.7, -5.8},
  {-1.5, -0.6, -5.9},
  {-1.4, -0.5, -6},
  {-1.6, -1, -6.5},
  {-1.4, -1, -6.4},
  {-1.2, -0.9, -6.8},
  {1.4, -0.6, -6.5},
  {4.5, -0.4, -5.5},
  {6.3, 2.6, -2.1},
  {6.3, 3.9, 1.4},
  {6.4, 5.5, 4.5},
  {6.4, 6, 7.1},
  {6, 4.9, 6.5},
  {1.7, 2.4, 2.1},
  {0.1, 1, -0.2},
  {0, 0.4, -1.5},
  {-0.2, 0.2, -2.5},
  {-0.7, 0, -3.4},
  {-0.8, -0.2, -3.8},
  {-1, -0.2, -4.3},
  {-1.6, -0.2, -5},
  {-1.1, 0, -5.4},
  {-1.4, -0.2, -5.8},
  {-1.5, -0.4, -5.9},
  {-0.9, -0.6, -6.3},
  {-1.9, -0.4, -6.5},
  {-1.6, -0.6, -6.8},
  {-1.9, -1.2, -6.9},
  {-1.7, -1.3, -7.2},
  {-1.6, -1.1, -7.3},
  {0.6, -0.2, -6.9},
  {4, -1.1, -6},
  {4.8, 1.7, -2.2},
  {4.7, 4, 1.4},
  {5.7, 4.5, 4.1},
  {5.5, 5.1, 6.5},
  {5, 3.4, 5.8},
  {2.3, 1.5, 2.3},
  {0.5, 0.4, -0.1},
  {-0.3, -0.2, -1.5},
  {-0.3, -0.7, -2.9},
  {-0.4, -0.9, -3.4},
  {-0.6, -1.1, -3.8},
  {-0.9, -1, -4.4},
  {-1.9, -0.5, -5.1},
  {-1.7, -0.5, -5.6},
  {-1.6, -1, -5.8},
  {-1.1, -1.5, -5.9},
  {-1.4, -1.6, -6.2},
  {-1.9, -1.9, -6.3},
  {-1.3, -1.7, -6.8},
  {-1.4, -1.4, -6.8},
  {-1.4, -2, -7},
  {-0.6, -1.8, -7},
  {2.1, -1.1, -6.5},
  {5, -0.5, -5.8},
  {6.1, 2.8, -1},
  {6.5, 4.1, 1.3},
  {6.8, 4.8, 4.8},
  {5.6, 4.7, 6.6},
  {4.4, 4.1, 5.8},
  {2.2, 1.9, 2.5},
  {1.4, 0.9, 0},
  {1.1, 0.3, -1},
  {0, 0, -2},
  {-0.4, -0.4, -2.6},
  {-1, -1, -3.4},
  {-1.1, -1.2, -2.7},
  {-1.4, -1.4, -2.4},
  {-2.5, -1.5, -2.8},
  {-2, -1.7, -3.6},
  {-2.4, -2, -4.5},
  {-2.1, -2.1, -5.1},
  {-2.2, -2.3, -5.7},
  {-2.2, -2.1, -6.1},
  {-2.3, -2, -6.5},
  {-0.9, -2.5, -6.8},
  {-0.8, -2.1, -6.7},
  {0.9, -1.5, -6.4},
  {3, -0.8, -5.5},
  {4.5, 2.2, -2.4},
  {5.4, 3.5, 0.2},
  {5.7, 4.2, 3.7},
  {5.4, 3.3, 5},
  {5.1, 3.4, 4.7},
  {3.8, 2, 2.9},
  {3.2, 1.2, 0.7},
  {2.3, 0.7, -0.7},
  {2.3, 0.5, -1.3},
  {3, 0.3, -1.7},
  {3.3, 0.2, -2.4},
  {3.3, -0.2, -2.8},
  {3, 0, -3.1},
  {3.2, -0.1, -3.2},
  {2.8, 0, -3.7},
  {3.3, 0.2, -4},
  {3.3, 0, -4},
  {3.8, 0.6, -4.1},
  {4.3, 0.9, -4.2},
  {3.3, 1, -4.2},
  {1.7, 0.7, -4.2},
  {2.3, 0.8, -4.6},
  {3.2, 0.8, -4.1},
  {4, 2.7, -3.1},
  {5.2, 2.5, -0.8},
  {6.7, 4.2, 1.7},
  {7.6, 4.5, 5.4},
  {7.9, 5.7, 7.4},
  {6.9, 5.5, 7.2},
  {5.3, 3.5, 4.1},
  {2.6, 2.7, 1.8},
  {4.4, 1.9, 0.1},
  {2.5, 1.4, -0.7},
  {2.6, 0.8, -1.5},
  {3.9, 0.4, -1.9},
  {3.9, 0.6, -2.4},
  {3.7, 0.9, -2.7},
  {3.6, 1, -2.9},
  {3.6, 0.9, -2.6},
  {4.1, 0.3, -2.5},
  {4.5, 0.4, -2.3},
  {4.6, 0.4, -1.8},
  {4.6, 0.7, -2},
  {2.4, 0.5, -2},
  {2.7, -0.1, -2.2},
  {4, 0.1, -1.8},
  {5.2, 0.5, -1.7},
  {5.5, 0.8, -0.8},
  {6.3, 0.9, 0.1},
  {7.2, 1, 1.4},
  {6.1, 1.4, 2.5},
  {6.2, 2, 3.5},
  {6.2, 1.3, 4.3},
  {6.5, 1.5, 3.1},
  {4.7, 1.6, 2.1},
  {3.3, 0.7, 1.8},
  {4.1, 0.9, 1.7},
  {4.4, 0.3, 1.5},
  {3.3, 1, 1.4},
  {2.9, 1.2, 0.8},
  {2.3, 0.9, -0.2},
  {2.2, 1, -0.3},
  {2.1, 1.3, -0.4},
  {1.7, 1.3, -0.1},
  {1.6, 1.8, 0.2},
  {1.1, 2.2, 0.5},
  {0.4, 1.7, 0.3},
  {0.3, 1.6, 0.2},
  {-0.2, 1.3, 0},
  {-0.1, 1.4, -0.2},
  {0.6, 2, -0.3},
  {2.5, 1.2, -0.3},
  {4.1, 1.6, 0.1},
  {4.5, 4.1, 0.6},
  {6.6, 6.5, 2.6},
  {5.9, 7.5, 5},
  {5.4, 7.2, 6.7},
  {3.4, 5.7, 4.1},
  {2.5, 3.8, 1.8},
  {1.6, 2.9, 0.5},
  {1.2, 2.3, -0.6},
  {0.9, 2.3, -1.1},
  {-0.5, 1.9, -1.8},
  {-1.8, 1.3, -2.2},
  {-1.1, 0.9, -2.9},
  {-1, 0.6, -3.4},
  {-1.9, -0.1, -4.2},
  {-1.9, 0.1, -4.5},
  {-0.9, 2.1, -4.7},
  {-0.1, 2.7, -4.7},
  {2.1, 2.6, -4.9},
  {2.1, 2.2, -5.2},
  {2.5, 2.1, -5.6},
  {1.7, 1.2, -6},
  {1.8, 2.1, -6},
  {4.9, 3.6, -5.1},
  {6, 5.6, -1.6},
  {6.2, 6.8, 1.5},
  {6.6, 7.6, 4.5},
  {6.5, 8, 6.3},
  {6.7, 7.6, 6.9},
  {2.5, 5.5, 4.4},
  {0.9, 4.1, 1.5},
  {0.6, 3.7, -0.3},
  {1.2, 3.5, -1.2},
  {0.9, 2.4, -2.3},
  {0, 1.8, -2.7},
  {0, 1.6, -3.3},
  {0.2, 1.7, -3.7},
  {0.6, 1.7, -3.7},
  {1.4, 2.1, -3.3},
  {0.6, 2, -2.7},
  {0.3, 1.3, -2.8},
  {0.1, 1.4, -3.2},
  {0.2, 1.5, -2.8},
  {0.4, 1.3, -2.8},
  {0.6, 0.9, -2.8},
  {1.4, 1.4, -2.7},
  {2, 1.3, -2.2},
  {2.6, 1.7, -1.2},
  {2.8, 2.1, -0.1},
  {3.2, 2.2, 0.7},
  {3, 2.1, 1.6},
  {3.6, 2.8, 3.4},
  {2.6, 2.2, 4.4},
  {1.3, 1.9, 2.8},
  {1.1, 1.6, 1.2},
  {0.9, 1.1, 0.1},
  {-0.2, 1.1, -0.8},
  {-1.1, 1.1, -1.7},
  {-0.3, 1.1, -1.8},
  {-0.2, 0.5, -1.8},
  {-1.2, 1.2, -1.8},
  {-0.8, 0.6, -2.2},
  {-1.4, 0, -3.3},
  {-1.1, -0.6, -3.3},
  {-1.2, -0.5, -3.7},
  {-1.1, 0.2, -4.3},
  {-1.2, -0.5, -5},
  {-1, -1.2, -5.1},
  {-1.5, -1.9, -5.4},
  {-0.9, -0.9, -5.8},
  {1.8, -1.2, -5.4},
  {5.4, 0, -4.7},
  {6.7, 2.6, -0.3},
  {7.8, 4.9, 2.6},
  {8.6, 6.6, 5.7},
  {8.3, 7.4, 8},
  {7.6, 6.2, 7.6},
  {3.7, 4.3, 3.9},
  {1.8, 3.1, 1.2},
  {2.2, 2.6, -0.1},
  {3.3, 3.3, -0.3},
  {2.9, 3.5, -0.3},
  {3.2, 3.7, -0.7},
  {2.5, 3.4, -0.7},
  {2.7, 2.8, -0.9},
  {1.5, 3, -0.9},
  {2, 2.4, -1},
  {2.4, 2, -0.9},
  {2.2, 2.2, -1},
  {0.9, 2.9, -1.1},
  {0.6, 2.3, -1.8},
  {0.2, 1.5, -2.5},
  {0.2, 1.4, -3.2},
  {0.1, 1.5, -3},
  {3.4, 1.7, -2.6},
  {6, 1.9, -2},
  {6.8, 4.3, 1.5},
  {6.9, 6.4, 5.1},
  {7, 7.5, 8.1},
  {7.1, 7.8, 10.2},
  {6, 6.3, 9.7},
  {4.3, 4.8, 6.2},
  {3.3, 3.5, 3.4},
  {3.2, 2.4, 1.1},
  {2.5, 2.4, 0},
  {2.5, 2.5, -0.6},
  {2.1, 2.4, -1},
  {2.3, 2.2, -1},
  {2.2, 2.5, -0.8},
  {2.4, 2.3, -1.4},
  {2, 2.2, -1.7},
  {1.6, 2, -1.5},
  {1.6, 1.5, -1.6},
  {1.7, 1.2, -1.1},
  {2, 0.8, -1.6},
  {1.7, 1.2, -2.1},
  {0.8, 1.6, -2},
  {1.1, 1.6, -1.4},
  {2.7, 1.9, -1.1},
  {4.7, 2.7, -0.9},
  {5.3, 4.3, 0.9},
  {6.9, 4.9, 3.7},
  {7.7, 5.6, 6.4},
  {7.1, 6.8, 8.7},
  {6.8, 5.8, 9},
  {4.9, 4.4, 5.2},
  {3.2, 3.7, 2.4},
  {1.7, 2.5, 0.8},
  {1.2, 2.1, 0},
  {2.4, 1.9, -0.6},
  {2.8, 2.7, -1.1},
  {2.9, 2.7, -0.7},
  {2.7, 2.6, -0.1},
  {2, 2.7, 0.3},
  {2.2, 2.7, 0.5},
  {1.3, 3, 0.3},
  {1.4, 2.7, 0},
  {1.8, 2.4, -0.4},
  {2, 2.4, -0.4},
  {2, 2.6, 0.2},
  {1.9, 2.8, 0.4},
  {2, 2.5, 0.7},
  {2.1, 2.8, 1},
  {2.1, 2.9, 1.1},
  {2.4, 3.3, 1.6},
  {2.4, 3.4, 2.7},
  {2.6, 3.7, 3.4},
  {3, 3.7, 4.3},
  {3, 3.9, 4.9},
  {2.7, 3, 4.5},
  {2.8, 2.2, 3},
  {2.8, 1.7, 1.5},
  {1.6, 1.6, 0.5},
  {1.1, 1.6, -0.3},
  {1, 1.4, -1.2},
  {1.3, 1.6, -1.4},
  {1.3, 1.9, -0.8},
  {1.5, 1.7, -1},
  {1.6, 1.6, -0.9},
  {1.4, 1.6, -1},
  {1.1, 1.6, -1.3},
  {0.5, 2.1, -1.6},
  {0.2, 2, -2.3},
  {0.3, 1.5, -2.6},
  {0.5, 1.3, -2.9},
  {0.7, 1.4, -2.8},
  {2.2, 2, -2.1},
  {3.5, 3.5, -0.9},
  {5.6, 5.9, 0.4},
  {6.7, 6.7, 3.3},
  {7.7, 7.9, 6},
  {7.3, 7.6, 8.1},
  {6.3, 7.4, 8.5},
  {4.5, 5.2, 7.1},
  {3.1, 4.5, 4.2},
  {2.4, 3.9, 2.8},
  {2.5, 3.6, 1.8},
  {2.6, 3.5, 1},
  {2.2, 3.6, 0.5},
  {2.4, 3.6, 0},
  {2.7, 3.3, 0},
  {1.6, 2.8, -0.7},
  {2.1, 2.3, -0.9},
  {1.6, 2.2, -1.6},
  {1.5, 1.9, -1.9},
  {2.3, 1.7, -2},
  {2.5, 1.6, -2.3},
  {2.9, 1.5, -2.3},
  {2.9, 1.3, -2.6},
  {3.2, 1.5, -2.8},
  {3.9, 2.1, -2.7},
  {4.1, 2.7, -1.6},
  {4.2, 3.3, -0.3},
  {4.7, 3.9, 0.9},
  {5.4, 4.6, 2.4},
  {6, 5.1, 3.7},
  {5.9, 4.7, 4.8},
  {5.2, 4.6, 4.7},
  {5.2, 4.5, 4.1},
  {4.8, 4.4, 3.5},
  {4.7, 4.3, 3.3},
  {4.4, 4.2, 3},
  {3.5, 4.2, 2.8},
  {3.6, 4, 2.8},
  {3.8, 3.7, 2.7},
  {4.7, 3.9, 2.7},
  {4.7, 3.8, 2.8},
  {4.7, 3.8, 2.9},
  {4.4, 3.9, 2.7},
  {4.6, 3.9, 2.7},
  {4.3, 3.2, 2.6},
  {4.3, 2.6, 2.6},
  {4.7, 2.7, 2.3},
  {5, 3, 0.9},
  {5.7, 3.5, 0.4},
  {7.7, 3.5, 0.7},
  {8.6, 5.9, 4.2},
  {8.7, 8, 7.5},
  {8.9, 9, 9.8},
  {7.2, 9.8, 11.7},
  {6.8, 8.7, 11.3},
  {6, 7.1, 9.3},
  {5.3, 6.2, 7},
  {5.1, 5.4, 5.4},
  {4.7, 5.6, 3.5},
  {4.4, 5.6, 3.6},
  {4.4, 5.7, 3.5},
  {4.4, 5.3, 3.8},
  {4.5, 5.1, 3.8},
  {4.4, 4.7, 3.7},
  {4.1, 4.4, 3.7},
  {3.7, 4.3, 3.7},
  {2.4, 4.5, 3.8},
  {1.8, 3.8, 3.9},
  {2, 3.8, 3.4},
  {5.5, 4.1, 2.8},
  {6.7, 4.5, 2.1},
  {4.9, 7, 1.9},
  {7.1, 8.2, 2.8},
  {10.8, 8.4, 5.4},
  {11, 9.2, 11.7},
  {11.9, 11.9, 14.9},
  {12.5, 13.7, 16},
  {12.7, 13.8, 16.6},
  {13.5, 13.7, 16.1},
  {8.9, 12.6, 11.7},
  {6.9, 10.8, 7.6},
  {7.2, 10, 5.5},
  {6.7, 9.6, 3.9},
  {5.7, 9.1, 2.9},
  {5.4, 7.8, 1.9},
  {5.3, 6.9, 1.4},
  {4.8, 7.1, 0.9},
  {4.6, 6.4, 0.1},
  {4.6, 6.4, 0.1},
  {4.6, 6, -0.5},
  {4.3, 5.7, -0.7},
  {4.5, 5.7, -1.1},
  {3.9, 5.3, -1.3},
  {4.3, 4.5, -1.7},
  {4.7, 4.6, -2},
  {5.5, 4.5, -1.9},
  {7.7, 5.7, -1.5},
  {11.1, 6, 0},
  {11.8, 7.2, 4.3},
  {12.5, 9.8, 8},
  {11.8, 10.8, 11.2},
  {12, 12.1, 13.1},
  {11.4, 11.3, 12.8},
  {7.9, 8.9, 8.8},
  {5.5, 7.1, 4.9},
  {4.7, 6, 2.7},
  {4.7, 5.4, 1.5},
  {4.1, 4.9, 0.9},
  {3.6, 4.2, 0},
  {3.5, 3.8, -0.4},
  {2.6, 3.5, -1.1},
  {1.6, 2.9, -1.4},
  {2.6, 2.6, -1.8},
  {1.2, 2.4, -2},
  {0.9, 2.1, -2.3},
  {0.9, 1.6, -2.6},
  {0.5, 1.7, -2.8},
  {1, 1.9, -2.8},
  {1.2, 2.2, -2.5},
  {2.2, 2.9, -2.6},
  {4.1, 2.7, -2.4},
  {7.2, 3.5, -1.3},
  {8.7, 4.3, 1.8},
  {9.6, 6, 5.1},
  {10, 7, 8},
  {9.9, 7.9, 10.2},
  {9.3, 8.3, 11.4},
  {6.6, 6.9, 7.6},
  {5.2, 5.8, 3.4},
  {4.7, 5.2, 1.6},
  {4.8, 5.4, 1},
  {4.5, 5.3, 0.1},
  {4.8, 5.2, -0.6},
  {5.9, 5.2, -1.1},
  {5.5, 5.3, -1.4},
  {5.1, 5, -1.6},
  {3.1, 5, -1.8},
  {4.2, 4.9, -2.3},
  {5.4, 4.4, -2.6},
  {4.9, 4.2, -2.9},
  {3.9, 3.6, -3},
  {3.6, 3.4, -3.2},
  {3, 3.1, -3.2},
  {3.1, 3.1, -3.5},
  {4.9, 3.3, -3.4},
  {8.5, 4, -1.8},
  {10, 6.3, 1.1},
  {10.7, 8.5, 4.8},
  {11.2, 8.9, 8.1},
  {10.7, 9.4, 10.9},
  {10, 9, 11.8},
  {7.1, 6.9, 7},
  {5.1, 5.7, 3.6},
  {4, 4.8, 2.1},
  {3.3, 4.4, 0.6},
  {3.2, 3.9, 0.2},
  {2.6, 3.7, -0.4},
  {2.3, 3.7, -1},
  {2, 3.8, -1.3},
  {2.3, 3.5, -1.6},
  {1.8, 3.1, -2.1},
  {2.1, 3.4, -2.2},
  {2.3, 3.7, -2.3},
  {1.5, 3.3, -2.4},
  {1.3, 3, -2.4},
  {1.2, 2.6, -2.7},
  {0.9, 2.1, -3.1},
  {1.5, 2.3, -2.9},
  {3.8, 2.4, -2.8},
  {5.9, 2.8, -2},
  {6.5, 6, 1.3},
  {6.3, 6.4, 1.9},
  {7.1, 6.9, 6.2},
  {7.1, 7.3, 8.5},
  {5.9, 6.7, 10.1},
  {4.6, 4.5, 6.8},
  {3.7, 3.8, 3.8},
  {3.4, 3.5, 2.2},
  {2.4, 2.9, 1.1},
  {2.3, 2.8, 0.2},
  {1.5, 2, 0},
  {0.6, 1.4, 0},
  {1.3, 1.1, -0.3},
  {1.8, 0.9, -0.4},
  {1.2, 1.5, -0.5},
  {1.1, 1.2, -0.7},
  {1.1, 1, -1.2},
  {1.3, 0.6, -1.8},
  {1, 0.6, -2.1},
  {0.1, 0.7, -2.4},
  {0.9, 0.7, -2.8},
  {1.2, 0.7, -3.2},
  {2.1, 1.5, -3},
  {2.9, 3, -1.9},
  {3.9, 2.9, -0.4},
  {4.8, 3.7, 1.1},
  {6.3, 5.6, 3.7},
  {6.1, 6.7, 6.8},
  {6.4, 6.9, 8.7},
  {4.1, 4.7, 6},
  {2, 3.4, 2.8},
  {1.5, 2.7, 1.1},
  {1.4, 2, 0.5},
  {1.3, 1.5, -0.4},
  {1.6, 1.3, -0.8},
  {1.8, 1.9, -1.2},
  {1.7, 2.1, -1.7},
  {1.4, 2, -1.7},
  {1.9, 1.7, -1.3},
  {1.2, 1.7, -0.7},
  {0.7, 2, -0.3},
  {1, 2.2, -0.3},
  {0.6, 1.7, -0.4},
  {0.4, 1.4, -0.7},
  {1.1, 1, -1.5},
  {3.7, 1.1, -1.8},
  {3.5, 1.8, -1.8},
  {5.1, 2.5, -0.6},
  {4.9, 2.8, 1},
  {4.8, 3.6, 1.9},
  {5.8, 3.5, 3.3},
  {6.5, 3, 4.9},
  {6.6, 3.5, 5.7},
  {5.1, 3.4, 5.5},
  {4.3, 3, 3.4},
  {5.1, 3, 1.9},
  {4.6, 2.9, 1.4},
  {4.5, 3.1, 1},
  {3.9, 3, 1.2},
  {4.2, 2.7, 0.9},
  {4.4, 2.8, 0.4},
  {4.6, 2.9, -0.1},
  {3.1, 2.6, -0.8},
  {2.7, 3, -1.3},
  {1.8, 2.4, -1.3},
  {2.9, 2.5, -1.3},
  {3.5, 2.2, -1.4},
  {5.1, 3.2, -1.2},
  {5.7, 4.6, -1.1},
  {7, 3.2, -0.8},
  {9.5, 6.1, -0.7},
  {11.9, 7.4, -0.1},
  {13.9, 8.4, 2.1},
  {15, 13, 5.7},
  {14.1, 15.6, 10.1},
  {15.5, 15.9, 12.9},
  {15.3, 17, 15.2},
  {14.4, 17, 15.4},
  {13.7, 17.3, 15.4},
  {12.7, 17.6, 14.2},
  {12.5, 17.4, 12.2},
  {11.1, 16.5, 10.2},
  {10.4, 14, 7.1},
  {10.9, 12.8, 5.7},
  {11.5, 12.4, 5},
  {10.7, 11.5, 3.3},
  {10.1, 11.6, 3.4},
  {9.9, 11.4, 2.6},
  {9.3, 11.2, 2.3},
  {8.8, 10.1, 2.1},
  {9.3, 10.5, 1.5},
  {8.6, 10.1, 1},
  {8.9, 9.7, 0.8},
  {9.8, 10, 1},
  {11.7, 11.3, 1.7},
  {12.7, 11.1, 3.4},
  {13.4, 11.1, 5.2},
  {14, 12.1, 7.7},
  {13.1, 12.5, 10},
  {12.8, 12.9, 12.9},
  {12.6, 12.4, 14.5},
  {9.2, 10.5, 11.8},
  {6.5, 8.9, 7.6},
  {5.7, 8, 5.1},
  {5.7, 7, 3.2},
  {4.1, 6.2, 2},
  {3.6, 5.1, 1.2},
  {2.7, 4.4, 0.9},
  {3.7, 4, 0.3},
  {4.8, 3.7, 0.9},
  {4.7, 3.5, 1.5},
  {5.1, 3.3, 1.8},
  {5.3, 3.6, 1.9},
  {4.9, 4.2, 1.8},
  {4.9, 4.1, 1.6},
  {4.8, 3.9, 1.6},
  {4.7, 3.9, 1.6},
  {4.7, 3.8, 1.8},
  {4.9, 4.3, 1.9},
  {5.3, 4.8, 2.5},
  {6.2, 4.8, 3.4},
  {7.2, 5.5, 4.6},
  {8.1, 7.3, 5.8},
  {8.3, 7.1, 7},
  {7.1, 7.2, 9.2},
  {5.9, 7, 9},
  {4.3, 5.9, 6.5},
  {3.2, 5.2, 4.3},
  {3.1, 5, 3},
  {2.8, 4.5, 3},
  {2, 4, 1.7},
  {3, 3.9, 1.4},
  {2.9, 3.9, 1.5},
  {3.6, 3.8, 1.4},
  {3.9, 4, 1.8},
  {4, 3.8, 2},
  {4.2, 3.6, 2.3},
  {4.8, 3.8, 2.4},
  {4.6, 3.8, 2.5},
  {4.1, 3.7, 2.4},
  {4.5, 4, 2.7},
  {4.5, 3.9, 2.6},
  {4.4, 3.9, 2.6},
  {4.6, 4.2, 3.2},
  {4.7, 3.9, 3.7},
  {5.1, 3.5, 3.9},
  {5.2, 3.2, 4},
  {5.9, 3.4, 4.6},
  {6.1, 3.3, 5},
  {5.2, 3.3, 5.2},
  {5, 3.3, 4.9},
  {4.6, 2.9, 4.4},
  {4.1, 2.9, 4.3},
  {3.9, 2.9, 4.1},
  {3.8, 3.2, 4},
  {3.8, 3.4, 4},
  {4.5, 3, 3.9},
  {5.7, 3.3, 3.9},
  {5.2, 3, 3.9},
  {4.1, 2.7, 3.9},
  {4.1, 2.6, 3.8},
  {4, 2.3, 3.8},
  {4.1, 2.4, 3.6},
  {4.1, 2.2, 3.3},
  {3.7, 1.9, 3.2},
  {3.9, 1.7, 3},
  {4.3, 2.1, 3},
  {4, 2.3, 3},
  {3.5, 2.2, 3},
  {2.5, 2.1, 3},
  {2.9, 2.1, 2.9},
  {3.1, 1.5, 2.7},
  {4.9, 1.2, 2.2},
  {5.8, 1.7, 2.1},
  {5, 1.9, 2},
  {5.2, 1.8, 2},
  {4.9, 1.7, 2.1},
  {4.5, 1.7, 2.2},
  {3.5, 1.9, 2.2},
  {3.2, 2.3, 2.2},
  {2.5, 2.4, 2.2},
  {1.3, 2.1, 2.2},
  {1.2, 2.3, 2.9},
  {0.9, 2.2, 3.5},
  {0.1, 1.7, 3.9},
  {-0.5, 1.3, 2.5},
  {-0.8, 0, 0.9},
  {0.2, 0, 0},
  {0.2, 0.4, -0.1},
  {0.2, 0.6, 0.3},
  {0.1, 1.4, 0.3},
  {0.9, 2.3, 1},
  {0.4, 2.9, 2.5},
  {1.1, 3.2, 3.6},
  {1.1, 2.7, 4.3},
  {0.5, 1.9, 4},
  {-0.1, 1.8, 4.8},
  {-0.5, 1.6, 4.1},
  {-1.3, 1, 2.7},
  {-1.5, 0.5, 2.3},
  {-2.1, 0, 1.7},
  {-3.4, -0.4, 2.1},
  {-3.8, -0.9, 2},
  {-4.6, -1.2, 1.1},
  {-4.7, -1.4, 1.1},
  {-4.4, -1.6, 0.7},
  {-4.8, -1.8, 0.9},
  {-4.9, -1.9, 0.9},
  {-5.2, -2.1, 0.1},
  {-4.7, -2.1, 0},
  {-4.6, -2.3, 0.1},
  {-4.4, -2.4, -0.3},
  {-4.2, -2.3, -0.5},
  {-3.6, -2.3, -0.6},
  {-3, -2, -0.1},
  {-2.5, -1.6, 1},
  {-2.1, -1, 1.9},
  {-1.1, -0.8, 2.5},
  {-1.4, -0.5, 2.7},
  {-1.2, -0.1, 3},
  {-2, 0, 3.3},
  {-2.3, 0, 3.3},
  {-2.8, -0.3, 2.6},
  {-3.3, -0.7, 1.9},
  {-3.5, -0.8, 1.3},
  {-3.7, -1.1, 0.8},
  {-3.5, -1, 0.5},
  {-3.5, -1.2, 0.5},
  {-3.2, -1.4, 0.2},
  {-3.4, -1.6, 0.2},
  {-3.6, -1.8, 0},
  {-3.8, -2, -0.1},
  {-4, -2.1, -0.2},
  {-4.2, -2.6, -0.6},
  {-4.1, -2.9, -1},
  {-4, -3.1, -1.1},
  {-4, -3, -1},
  {-3.9, -2.8, -1},
  {-3.7, -2.7, -0.9},
  {-3.8, -2.3, -0.7},
  {-3.4, -2.3, -0.7},
  {-3.4, -2.2, -0.6},
  {-3.2, -2, -0.2},
  {-3.1, -1.2, 0},
  {-3.5, -1.2, 0.4},
  {-3.6, -1.7, 0.3},
  {-3.9, -2.9, -0.7},
  {-5.8, -3.2, -1.7},
  {-6.1, -3.5, -2},
  {-6.3, -3.7, -2.9},
  {-6.9, -3.8, -3.6},
  {-7.2, -3.8, -4.1},
  {-7.2, -3.8, -4.4},
  {-7.5, -4.4, -4.5},
  {-7.4, -4.5, -4.7},
  {-7.7, -4.8, -5.5},
  {-7.6, -4.6, -5.7},
  {-8, -5.1, -6.1},
  {-8.4, -5.3, -6.6},
  {-8, -5.3, -6.9},
  {-8, -4.9, -7.3},
  {-7.6, -5.6, -7.2},
  {-4.3, -3.4, -7.1},
  {-0.6, -1.8, -5.8},
  {1.3, 0.8, -3.1},
  {2.8, 2.9, -0.8},
  {3.5, 3.9, 1.6},
  {3.5, 4.3, 4.2},
  {3.3, 4.6, 6.2},
  {1.9, 3.4, 6},
  {1.3, 2.4, 2.4},
  {0.3, 2.3, 1.3},
  {-1.2, 2.2, 0.4},
  {-1.7, 1.8, -0.2},
  {-1.8, 1.2, -0.6},
  {-2.2, 0.5, -1.7},
  {-1.9, 0.4, -2.3},
  {-2.4, 0.6, -3},
  {-2, 0.6, -3.7},
  {-2.4, 0.2, -3.8},
  {-2.3, -0.1, -4.4},
  {-2.4, -0.3, -4.6},
  {-2.7, -1, -4.8},
  {-2.8, -0.8, -5.1},
  {-2.3, -0.4, -5.3},
  {-0.9, -0.6, -5.1},
  {1.5, -0.9, -4.3},
  {3.3, -0.2, -1.8},
  {4.4, 3.9, 0.8},
  {5.2, 3.8, 3.3},
  {5.7, 5.3, 6.4},
  {5.7, 6.1, 8},
  {5.4, 7, 9.1},
  {3.3, 5.7, 6.4},
  {0.6, 2.7, 2.9},
  {0.7, 1.1, 0.9},
  {0.3, 0.5, 0.2},
  {-0.6, 0, -0.7},
  {-0.5, 0, -1.5},
  {-0.6, -0.5, -1.8},
  {-0.8, -0.8, -2.3},
  {-1.5, -1, -2.7},
  {-1.8, -1, -2.9},
  {-1.8, -0.6, -3.2},
  {-1.5, -0.6, -3.7},
  {-1.1, -1.1, -4.1},
  {-0.9, -0.2, -4.4},
  {-0.1, -0.6, -4.6},
  {0.5, -0.1, -4.8},
  {1.1, 0.1, -4.7},
  {3.2, -0.3, -4.1},
  {5.4, -0.4, -3.1},
  {7.7, 3.9, -1.5},
  {8.5, 7.2, 0.6},
  {10, 9.8, 2.6},
  {10.5, 9, 5.9},
  {11, 11.4, 8.6},
  {7.4, 9.7, 6.7},
  {4, 7.2, 2.9},
  {3.8, 6.5, 1.3},
  {3.3, 6, 0.3},
  {3.6, 5.1, -0.2},
  {2.9, 4.6, -0.7},
  {3, 3.7, -1.2},
  {2, 3.8, -1.8},
  {1.7, 3, -2.4},
  {1.3, 2.3, -2.7},
  {0.8, 2.3, -3},
  {0.3, 2.1, -3.4},
  {0.2, 1.7, -3.8},
  {-0.4, 1.2, -4.1},
  {-0.4, 1.1, -4.2},
  {-0.5, 1.5, -4.6},
  {0, 1.6, -4.6},
  {3.1, 2.1, -4.6},
  {6.3, 2.6, -2.8},
  {7.6, 6.9, 1.3},
  {7.1, 7.5, 4.8},
  {8, 6.7, 8.2},
  {8.5, 8.7, 10.4},
  {7.8, 8.6, 11.5},
  {5.8, 7.3, 8.6},
  {2.5, 4.5, 4.1},
  {1.8, 3.2, 2},
  {1.8, 3.2, 0.6},
  {1.7, 2.3, -0.1},
  {1.2, 2.4, -0.8},
  {1.2, 2.3, -1.4},
  {1.6, 2, -1.8},
  {0.6, 2.1, -2.1},
  {0, 1.7, -2.6},
  {-0.1, 1.1, -2.7},
  {-0.7, 0.5, -3.2},
  {-1.1, 0.2, -3.5},
  {-0.6, -0.1, -3.9},
  {-0.4, -0.1, -4.3},
  {-0.8, -0.1, -4.5},
  {-0.2, 0, -4.4},
  {2.8, 0.5, -4.4},
  {5.2, 3.5, -3},
  {6, 4.2, 1.3},
  {6.5, 5.8, 4.2},
  {7.1, 7, 7.7},
  {7.4, 7.7, 9.6},
  {6.4, 7.7, 10},
  {4.4, 5.9, 8},
  {2.5, 3.3, 4.2},
  {1.2, 2.8, 2.9},
  {0, 1.5, 1.2},
  {-0.6, 1.3, 0},
  {-0.6, 1.1, -0.9},
  {-0.7, 0.8, -1.4},
  {-0.4, 0.7, -1.9},
  {-0.8, 0.2, -2.3},
  {-0.5, 0.3, -2.6},
  {-1.3, 0.5, -2.5},
  {-0.6, 0.6, -3},
  {-0.5, -0.2, -3.1},
  {-0.2, 0.2, -3.7},
  {-0.5, 0.5, -3.9},
  {0.6, -0.5, -4.1},
  {2, -0.5, -3.9},
  {5.6, 0.3, -3.5},
  {7.9, 2, -2.2},
  {10, 4.4, 0.7},
  {10.2, 5.9, 3.9},
  {10.9, 7.6, 6.7},
  {10.9, 8.5, 8.2},
  {10, 9.4, 7.9},
  {6.5, 7.8, 5.3},
  {4.8, 5.1, 2.9},
  {2.4, 4, 1.8},
  {4.2, 4.4, 0.7},
  {5.3, 4.5, 0.1},
  {4.9, 4.7, -0.5},
  {4.2, 4.3, -0.9},
  {3.7, 3.6, -1.2},
  {4.1, 2.9, -1.6},
  {3.8, 2.7, -1.7},
  {4.1, 2.8, -1.5},
  {3.9, 2.9, -1.3},
  {3, 2.7, -1.2},
  {1.3, 2.4, -1.3},
  {1, 1.6, -1.8},
  {0.6, 1.5, -2},
  {1.2, 1.8, -2.7},
  {4.5, 2.1, -2.7},
  {6.9, 3.1, -1.1},
  {7.8, 6.9, 2.1},
  {8.5, 7.9, 6.3},
  {9.3, 9.4, 9.9},
  {9.5, 10.2, 12.3},
  {9.1, 10.5, 13.8},
  {6.8, 9.1, 11.1},
  {4, 6.3, 6.7},
  {3, 4.8, 3.3},
  {1.9, 3.9, 2},
  {1.6, 3.3, 1.1},
  {1.4, 3, 0.2},
  {1.4, 3.5, -0.4},
  {1.4, 3.3, -0.7},
  {1.3, 2.9, -1.3},
  {1.6, 2.1, -1.6},
  {2, 2.1, -1.7},
  {2.8, 1.9, -2.1},
  {2.9, 2.1, -2.3},
  {2.5, 2.7, -2.5},
  {3.3, 2.3, -2.7},
  {3.4, 2.5, -2.9},
  {4.1, 1.7, -3.2},
  {7.9, 2.8, -2.6},
  {10.2, 4.7, -1.2},
  {11.6, 10.7, 2.9},
  {12.2, 11.8, 6.8},
  {12.6, 12.7, 10.6},
  {12.7, 13.3, 14},
  {12.2, 13, 16.2},
  {10.9, 11.4, 14.2},
  {8.2, 9.8, 9.9},
  {6.8, 9.3, 8},
  {6.9, 9, 5.3},
  {6.6, 8, 3},
  {5.3, 6.9, 2.1},
  {3.9, 6.2, 0.6},
  {3.8, 5.5, 0.1},
  {2.2, 5.3, -0.4},
  {1.5, 4.7, -1},
  {1.9, 3.6, -1.6},
  {2.3, 2.9, -2},
  {1.3, 1.9, -2.7},
  {0.9, 1.1, -2.9},
  {0, 1, -3.5},
  {-0.2, 0.3, -3.4},
  {-0.5, 0.9, -3.5},
  {2.1, 1.5, -3.6},
  {3.9, 3, -1.6},
  {4.5, 4.7, 1.7},
  {5.6, 6.1, 4.5},
  {6.2, 7.1, 7.6},
  {6.4, 8, 10.4},
  {6.5, 8.2, 10.4},
  {4.8, 7, 8.6},
  {1.4, 4, 5.1},
  {0.7, 2.9, 2.2},
  {0.8, 2.2, 0.6},
  {0.1, 1.7, -0.3},
  {-0.3, 1.4, -1},
  {-0.6, 1.1, -1.7},
  {-0.1, 1.1, -2.2},
  {0.3, 0.4, -2.5},
  {0.1, 0.2, -3.1},
  {-0.4, 0.2, -3.6},
  {-1, 0.3, -4.1},
  {-0.8, 0.4, -4.1},
  {-0.8, 0, -4.6},
  {-0.7, -0.6, -4.9},
  {-0.9, -0.8, -5},
  {0, -0.1, -5},
  {3.4, -0.3, -4.7},
  {5.8, 0.9, -2},
  {6.4, 4.1, 0.8},
  {7.1, 5.2, 4.5},
  {7.2, 6.7, 7.6},
  {7.2, 7.5, 10.4},
  {6.8, 7.5, 10.4},
  {5.8, 6.7, 7.7},
  {3, 4.4, 5.5},
  {1.8, 3.1, 2.7},
  {1.6, 2.7, 1.4},
  {1.5, 1.9, 0.5},
  {1.3, 1.4, -0.1},
  {0.1, 1, -0.9},
  {0.3, 0.6, -1.6},
  {1.8, 0.3, -2},
  {1.8, 0.1, -2.3},
  {2, 0.6, -2.9},
  {1.8, 0.4, -3.2},
  {1.3, 0.2, -3.5},
  {1.9, 0.5, -3.2},
  {2.5, 0.1, -2.4},
  {3.6, 0, -2.1},
  {3.8, 0, -2.6},
  {2.7, 0.1, -2.2},
  {2.6, 0.6, -0.8},
  {2.3, 1.8, 0},
  {2.1, 3, 1.9},
  {2.1, 3.6, 3.3},
  {2.1, 3.6, 4.8},
  {1.9, 3.6, 4.7},
  {1.7, 3.7, 4.8},
  {1.3, 3.4, 4.1},
  {1.2, 3.3, 3.5},
  {1.3, 3.1, 3},
  {1.3, 2.8, 2.7},
  {1.2, 2.4, 2.4},
  {1.2, 2.3, 2.3},
  {1.2, 2.2, 2.3},
  {1.2, 2, 2.2},
  {1.2, 1.6, 2.2},
  {1.1, 1.7, 2.2},
  {1.1, 1.7, 2.1},
  {0.9, 1.6, 2},
  {0.8, 1.6, 2},
  {0.1, 1.3, 2.1},
  {-0.2, 1.2, 2.1},
  {-0.2, 1.5, 2.2},
  {0.4, 2.1, 2.6},
  {0.9, 3.2, 3.1},
  {1.6, 3.3, 4.2},
  {2.4, 4, 5.9},
  {3.1, 4.4, 6.9},
  {3.7, 4.8, 7.3},
  {4.2, 4.7, 6},
  {3, 4.3, 5.5},
  {1.5, 3.8, 5.2},
  {1.8, 3.4, 4.7},
  {1.5, 2.9, 4.6},
  {1.6, 3.4, 4.6},
  {1.6, 3.2, 4.4},
  {1.5, 3.1, 4.1},
  {1.4, 3, 4.1},
  {1.3, 2.7, 3.7},
  {1.6, 2.7, 3.9},
  {1.6, 2.6, 3.7},
  {1.7, 2.5, 3.5},
  {1.6, 2.5, 3.4},
  {1.5, 2.4, 3.4},
  {1.5, 2.4, 3.3},
  {1.5, 2.4, 3.2},
  {1.5, 2.4, 3.3},
  {1.7, 2.7, 3.6},
  {2.3, 3, 4},
  {2.5, 3.4, 4.4},
  {3.4, 3.7, 5.4},
  {4.3, 4.1, 5.9},
  {4.7, 4.4, 6.4},
  {4, 4.4, 6.4},
  {4, 4, 6},
  {3.6, 3.8, 5.9},
  {3.1, 3.5, 5.3},
  {2.6, 3.6, 5.1},
  {2.3, 3.4, 4.9},
  {1.8, 3.1, 4.6},
  {1.1, 2.8, 4.2},
  {0.9, 2.7, 3.7},
  {1.1, 2.3, 3.5},
  {1.4, 2.1, 3.4},
  {1.6, 2.1, 3.2},
  {2, 2.1, 3},
  {1.8, 2.2, 2.9},
  {1.7, 2.3, 2.8},
  {1.4, 2.3, 2.8},
  {1.1, 2.2, 2.6},
  {0.7, 2.6, 1.7},
  {2, 2.8, 1.5},
  {2.9, 3.3, 2.2},
  {3.9, 4.7, 2.8},
  {4.5, 6.4, 4.8},
  {5, 7.3, 8.5},
  {6.1, 7.1, 10.5},
  {6.6, 7.7, 11.2},
  {5.8, 7.6, 10.6},
  {3.5, 4.4, 7.7},
  {2.5, 3.3, 5.1},
  {2.8, 3.1, 3.5},
  {2.8, 3.2, 3.1},
  {3.1, 3.6, 3.4},
  {1.7, 4, 3.2},
  {1.5, 4.1, 3.3},
  {0.8, 3.8, 3.2},
  {1.6, 3.3, 3},
  {1.6, 3.1, 2.5},
  {0.8, 2.8, 2.2},
  {1.6, 2.8, 2.2},
  {2, 3, 2},
  {1.8, 2.8, 1.9},
  {2.2, 2.8, 1.9},
  {2.5, 2.9, 2.2},
  {3.1, 3.7, 2.6},
  {3.5, 4.7, 3.7},
  {4.3, 5.5, 5.1},
  {5.4, 6.2, 6.9},
  {5.8, 6.9, 8.4},
  {6.1, 7.3, 10.5},
  {5.9, 6.8, 10.6},
  {4.8, 6.1, 10.4},
  {2.5, 5.6, 8.7},
  {1.6, 5, 7.5},
  {2.1, 4.7, 6.1},
  {1.8, 3.9, 4.6},
  {1.7, 3.5, 3.1},
  {1.9, 3.8, 2.4},
  {1.5, 4, 2.2},
  {1.7, 3.7, 1.9},
  {1.2, 3.6, 1.6},
  {0.4, 3, 0.7},
  {0.1, 2.6, 0.2},
  {-0.1, 2.3, -0.5},
  {0.2, 1.3, -0.7},
  {0.2, 0.7, -1.2},
  {0.6, 0.6, -1.5},
  {1.7, 1.2, -1.7},
  {4.1, 2.1, -1.2},
  {5.8, 3.6, 0.7},
  {5.8, 4.5, 2.8},
  {5.8, 4.7, 4.6},
  {6.9, 6.4, 6.6},
  {7.3, 8.1, 9.7},
  {7.8, 8.8, 10.5},
  {5.9, 8.1, 10.5},
  {4.4, 6.1, 8},
  {3.1, 4.9, 4.7},
  {1.8, 3.6, 2.6},
  {2.5, 2.9, 1.2},
  {1.4, 2.4, 0.5},
  {0.2, 2.1, -0.1},
  {0, 1.6, -0.6},
  {-0.1, 1.5, -1.1},
  {-0.6, 1.4, -1.4},
  {0.4, 1.4, -2},
  {0.9, 1.2, -1.9},
  {1.3, 1.7, -1.4},
  {1.3, 1.6, -1},
  {0, 1.3, -0.8},
  {0.8, 1.2, -1.3},
  {1.2, 1.8, -1.1},
  {4.3, 2.5, -1},
  {5.8, 3.3, 1.2},
  {5.6, 5.1, 3.7},
  {6.6, 6.3, 5.9},
  {6.7, 7.3, 7.4},
  {5.6, 6.6, 8.7},
  {4.3, 6.9, 9.4},
  {3.3, 6, 8},
  {2.8, 4.4, 7},
  {1.4, 3, 5.5},
  {0.8, 2.5, 4.6},
  {0.7, 2, 3.9},
  {0.5, 1.6, 3.5},
  {0.3, 1.2, 3.1},
  {0.3, 1.5, 2.9},
  {0.7, 1.8, 2.8},
  {0.9, 2.3, 2.5},
  {1.2, 3.3, 2.1},
  {1.5, 3.8, 1.8},
  {1.3, 4.3, 1.5},
  {1.3, 4.5, 1.1},
  {0.9, 3.1, 0.9},
  {0.7, 2.2, 0.3},
  {1, 2.7, 0.6},
  {3.3, 2.8, 1},
  {5.7, 4.6, 1.7},
  {7.8, 8.7, 2.4},
  {8.9, 10, 4.6},
  {9.8, 11.1, 8.7},
  {10, 11.9, 12.2},
  {10.3, 12.4, 13.9},
  {8.3, 11.2, 13.1},
  {4.7, 9, 8.4},
  {4.4, 9.5, 5.8},
  {3.8, 8.2, 3.6},
  {3.3, 6.5, 2.2},
  {2.5, 6.2, 1.1},
  {2.6, 5, 0.4},
  {2.4, 3.9, -0.4},
  {2.6, 3.8, -0.7},
  {1.4, 2.7, -1.3},
  {0.4, 2.8, -1.8},
  {-0.4, 2.6, -2},
  {-0.4, 1.8, -2.6},
  {0, 1.4, -2.9},
  {0.2, 0.9, -3},
  {0.9, 0.7, -3.5},
  {1.6, 1.2, -3.2},
  {3.9, 2.7, -2.5},
  {4.5, 4.6, -0.4},
  {6.6, 4.1, 1.3},
  {6.3, 4.1, 4.4},
  {6.7, 5.1, 6},
  {6.5, 5.7, 8},
  {5.7, 5.7, 8.7},
  {5.3, 5.2, 8.6},
  {4.1, 4.8, 7.8},
  {3.8, 4.6, 5.7},
  {3.3, 4.8, 4.7},
  {3.5, 4.4, 4},
  {3.4, 4.1, 3.4},
  {2.9, 3.9, 3},
  {2.4, 4, 2.6},
  {2.1, 4.1, 2},
  {2.6, 3.5, 1.3},
  {2, 3.3, 0.6},
  {1.8, 3, 0.3},
  {1.7, 2.7, -0.2},
  {1.9, 2.7, -0.4},
  {2, 2.7, -0.1},
  {2.3, 3, 0},
  {3.7, 4.3, 0.1},
  {4.7, 4.2, 0.8},
  {6.7, 7, 2.3},
  {8.3, 8.1, 6},
  {8.5, 9.1, 8.8},
  {9.6, 12.8, 10.6},
  {11.9, 13.8, 13.5},
  {11.4, 13.9, 15.7},
  {9.6, 12.5, 14.5},
  {6.5, 10.1, 10.2},
  {5.4, 9.2, 6.5},
  {4.2, 8.4, 4.1},
  {3.6, 7.6, 2.4},
  {3.2, 6.9, 1.4},
  {2.8, 6.9, 0.5},
  {2.6, 6, 0},
  {2.1, 5.3, -0.5},
  {2, 4.9, -1},
  {1.9, 4.5, -1.5},
  {1.4, 3.9, -1.9},
  {1.4, 3.2, -2.3},
  {1.3, 3.2, -2.7},
  {1.1, 2.3, -2.9},
  {1.2, 1.6, -3},
  {2.2, 1.9, -3.1},
  {6.8, 2.8, -3},
  {7.9, 5.4, 0.1},
  {8.1, 8.6, 4.7},
  {8.6, 10.3, 9},
  {9.4, 11.1, 12.2},
  {9.5, 11.9, 13.2},
  {8.8, 11.3, 12.5},
  {6.5, 9.6, 11.1},
  {4.9, 7, 9},
  {4.3, 5.8, 7.6},
  {3.5, 5.4, 4.9},
  {3.9, 4.2, 3.6},
  {3.1, 3.9, 3.9},
  {1.1, 5, 3.8},
  {1.1, 3.3, 2.4},
  {0.7, 2.5, 1.2},
  {0.2, 2.1, 0.2},
  {0.1, 2, -0.3},
  {-0.2, 1.6, -0.8},
  {-0.4, 1.3, -1.4},
  {-0.5, 1.5, -1.7},
  {0.6, 1.4, -1.9},
  {-0.1, 1, -2.4},
  {0.8, 1.5, -2.3},
  {3.9, 2.8, -1.2},
  {4.7, 4.7, 0.1},
  {4.2, 5.7, 0.5},
  {4.4, 6.2, 2.8},
  {5.1, 6.8, 6},
  {5.2, 7.3, 8.6},
  {5, 7.9, 8.9},
  {4.5, 7.3, 9},
  {2, 5.2, 7.6},
  {0.4, 4, 4},
  {1.6, 3.6, 2.1},
  {2.6, 3.2, 0.8},
  {2.7, 3.9, 1.2},
  {2.2, 4.5, 1.4},
  {2.2, 4, 1.7},
  {1.6, 3.5, 1.7},
  {0.6, 2, 1.1},
  {0.2, 1.3, -0.1},
  {-0.8, 1.3, -0.8},
  {-1.4, 0.7, -1.5},
  {-1.6, 0.3, -2},
  {-1.3, 0.2, -2.3},
  {-0.7, 0.1, -2.5},
  {0.3, 1, -2.8},
  {1.2, 2.4, -2.1},
  {1.7, 3.5, -0.2},
  {2.4, 4.7, 2},
  {4.6, 6.1, 6},
  {5.4, 7.1, 8.5},
  {5.7, 8.1, 9.6},
  {5.3, 8, 9.1},
  {3.2, 6.7, 7.9},
  {1.5, 4.4, 6},
  {1.1, 3.2, 4.6},
  {-0.4, 2, 1.5},
  {0.5, 1.5, 0.4},
  {0.3, 0.9, -0.6},
  {0.3, 0.4, -1.1},
  {0.2, 0.2, -2},
  {-1.3, 0, -2},
  {-2.1, -0.5, -2.4},
  {-2.3, -0.6, -2.8},
  {-2.7, -0.6, -2.9},
  {-2.8, -0.4, -3.5},
  {-2.8, -0.7, -4},
  {-3, -1.1, -4.3},
  {-2.9, -0.9, -4.4},
  {-1.9, -0.1, -4.1},
  {1.4, 0.6, -3.5},
  {3.5, 2, -0.7},
  {5.5, 3.5, 2.3},
  {5.7, 5.3, 6.3},
  {6.4, 7.1, 8.9},
  {6.7, 8.2, 10.2},
  {7.1, 9, 11.2},
  {6.4, 8.6, 10.1},
  {2.9, 6.2, 8},
  {1.6, 4.6, 4.6},
  {1.3, 3.4, 2.5},
  {0.6, 3, 0.8},
  {1.6, 2.2, -0.2},
  {1.7, 1.9, -0.7},
  {1.8, 1.4, -1.5},
  {1.8, 1.1, -1.8},
  {1.1, 1, -2.3},
  {0.6, 1.6, -2.6},
  {1.4, 1.5, -3.1},
  {1.2, 1, -3.1},
  {0.7, 0.6, -3.7},
  {0, 0.4, -3.9},
  {0, 0.2, -4.1},
  {0.8, 0.7, -4.2},
  {4.3, 2.2, -3.2},
  {5.2, 4.8, 0.1},
  {6.5, 6.8, 3.8},
  {8.3, 7.4, 8},
  {9.1, 9.1, 11.1},
  {9.5, 10.6, 13.2},
  {9.8, 11.4, 13.3},
  {8.7, 11.2, 12.5},
  {5.4, 8.7, 11},
  {3.4, 6.5, 6.8},
  {3, 5.8, 3.3},
  {2.3, 4.9, 1.6},
  {2.2, 3.8, 0.5},
  {4.5, 3.6, 0},
  {5.1, 4.4, -0.3},
  {4.7, 4.3, 0},
  {5, 4.2, 0.5},
  {4.8, 4, 0.6},
  {4.4, 3.9, 0.5},
  {2.7, 3.6, -0.3},
  {2.1, 3.1, -1.3},
  {1.8, 3.4, -1.9},
  {2.5, 3.9, -1.6},
  {3, 3.9, -1.4},
  {4.9, 5.2, 0.2},
  {6.9, 5.7, 3.4},
  {9.2, 6, 5.9},
  {11.1, 8.7, 10.3},
  {10.6, 10.6, 12.6},
  {9.9, 11.8, 14.3},
  {9.1, 11.6, 11.9},
  {7.8, 9.7, 11.1},
  {6.9, 8.8, 10.2},
  {4.9, 8.1, 9.4},
  {5.1, 7.5, 7.2},
  {4.3, 7.4, 5.1},
  {4.3, 6.6, 3.5},
  {3.3, 6, 3.2},
  {3.5, 6.5, 3},
  {3.7, 6.1, 2.8},
  {4, 5.7, 2.6},
  {4.3, 5.6, 3},
  {4.1, 5.1, 3.1},
  {3.3, 5.3, 2.9},
  {3.9, 5.4, 2.9},
  {4.1, 4.9, 2.5},
  {4.2, 5.1, 2.2},
  {4.9, 5, 3},
  {5.6, 6.2, 4.5},
  {5.9, 7.2, 6.6},
  {7.5, 8.5, 8.2},
  {9.2, 9.8, 9.5},
  {9.5, 10.9, 11.1},
  {9.1, 12, 13},
  {8.2, 11.9, 12.2},
  {6.8, 10.4, 11},
  {6, 8.7, 10},
  {4.9, 7.7, 8.7},
  {4.5, 7, 5.9},
  {3.5, 6.1, 5.4},
  {3.2, 5.4, 4.1},
  {2.7, 4.8, 2.4},
  {1.9, 4.8, 1.6},
  {2, 5.5, 1.2},
  {2.2, 5.6, 1.1},
  {2.6, 5.3, 1.9},
  {3.2, 5.3, 2.3},
  {3.9, 5.2, 2.8},
  {4.1, 5.6, 3.1},
  {4.2, 5.1, 3.3},
  {4.2, 5.3, 3.3},
  {4.5, 5.7, 3.5},
  {4.7, 6, 4},
  {5.6, 6.4, 4.6},
  {6.4, 7.9, 5.4},
  {7.3, 8.6, 7.4},
  {7.1, 8.8, 9.3},
  {7.7, 9, 10.8},
  {7.7, 8.9, 11.3},
  {6.7, 9.1, 11.3},
  {6, 8.2, 10},
  {4.9, 7, 9.1},
  {4.7, 7.3, 7.5},
  {4.1, 6.8, 6.8},
  {3.7, 6.7, 6.2},
  {3.9, 6.8, 5.7},
  {3.8, 6.7, 5.6},
  {4.4, 6.8, 5.5},
  {4, 6.2, 5.3},
  {3.3, 6.1, 4.7},
  {2.9, 5.9, 3.8},
  {2.9, 5.4, 3.7},
  {3, 5.1, 3},
  {3.5, 5.1, 2.7},
  {4.1, 5.6, 2.9},
  {4.8, 6.3, 3.4},
  {5.3, 6.4, 4.1},
  {5.1, 7.1, 5.2},
  {5.9, 7.7, 6.1},
  {5.8, 8.8, 8.1},
  {5.7, 9.2, 10.1},
  {5.7, 8.8, 9.8},
  {5.8, 8.6, 9.5},
  {6, 7.8, 9.3},
  {5.4, 7.4, 9.1},
  {4.4, 7.3, 8.6},
  {4.3, 7, 8.2},
  {4.2, 6.7, 7.7},
  {4.1, 6.5, 6.6},
  {4, 5.8, 5.1},
  {3.9, 5.7, 5.4},
  {3.6, 5.6, 5.3},
  {3.2, 5.4, 5},
  {3.3, 5.1, 4.3},
  {3.7, 4.8, 3.8},
  {3.6, 4.8, 3.7},
  {3.4, 4.8, 3.3},
  {3.1, 4.6, 2.6},
  {3.4, 4.7, 2.9},
  {3.9, 5, 3.2},
  {4.1, 4.9, 4.1},
  {4.9, 5.3, 5.4},
  {5.8, 5.8, 6.8},
  {6.2, 6.7, 7.8},
  {6, 7.6, 8.8},
  {5.4, 7.8, 9.4},
  {4.8, 6.9, 8.7},
  {4.4, 6, 8},
  {4, 5.5, 7.3},
  {3.7, 5.3, 6.8},
  {3.5, 5, 6.3},
  {3.3, 4.8, 6},
  {2.7, 4.5, 5.7},
  {2.6, 3.9, 5},
  {3, 3.7, 4.4},
  {3.3, 3.7, 4.4},
  {3, 3.3, 4.4},
  {2.3, 3, 4.2},
  {1.3, 2.7, 3.7},
  {0.5, 2.6, 2.7},
  {0.2, 2.5, 2.6},
  {0.2, 2.3, 2.6},
  {0.2, 2.3, 2.6},
  {0.9, 2.6, 2.8},
  {3.9, 3.1, 3.2},
  {5.9, 5.4, 3.7},
  {7.5, 6.6, 5.6},
  {8.5, 8.4, 8.1},
  {9, 9.8, 10.6},
  {9.5, 10.4, 12.8},
  {10.1, 10.5, 13.7},
  {8.5, 9.9, 13.4},
  {5.6, 7.9, 11.3},
  {3.4, 6.6, 9},
  {3.1, 6.1, 6.3},
  {2.9, 5.2, 4.2},
  {2.7, 4.7, 2.9},
  {2, 4.1, 1.8},
  {1.7, 4.3, 1.3},
  {1.8, 3.6, 0.6},
  {1, 3.3, 0.2},
  {1.5, 3.4, -0.3},
  {1.5, 2.9, -0.7},
  {0.5, 2.5, -1.1},
  {0.4, 3.4, -1.3},
  {0.7, 2.6, -1.8},
  {2.5, 2.4, -2.2},
  {3.4, 2.8, -2.1},
  {6.2, 4.2, -1.3},
  {7.7, 6.5, 2.4},
  {8.7, 8.8, 5.8},
  {9, 9.8, 9.8},
  {9.8, 10.8, 12.7},
  {10, 11.4, 13.5},
  {9.8, 11.5, 14.2},
  {9.2, 11, 12.8},
  {7.5, 9.7, 11.1},
  {5.5, 7.9, 10.6},
  {4.1, 8, 8},
  {3.1, 7.7, 5.7},
  {3.5, 6.9, 3.6},
  {3.5, 5.7, 2.5},
  {2.6, 4.7, 1.6},
  {2.4, 4.3, 0.8},
  {2.1, 4.1, 0.4},
  {2.1, 3.5, 0},
  {1.9, 3.2, -0.1},
  {1.4, 3.2, -0.4},
  {1.5, 3.1, -0.6},
  {0.9, 2.5, -1},
  {1.3, 3.3, -1.3},
  {3.2, 3.5, -1},
  {5.9, 3.8, 0.3},
  {6.7, 4.9, 4.2},
  {6.5, 5.8, 7.8},
  {6.5, 7.3, 9.6},
  {7.2, 8.2, 10.3},
  {9.2, 9.8, 10.8},
  {9.3, 10.7, 12.2},
  {8.3, 10.3, 11.8},
  {5.9, 9, 9.9},
  {3.4, 6.3, 7.1},
  {3.4, 5.6, 4.9},
  {4, 4.8, 3.4},
  {4.1, 4.5, 2.4},
  {4, 4.3, 3} ;
}
